* NMOS/PMOS models from
* https://people.rit.edu/lffeee/SPICE_Examples.pdf

.model EENMOS NMOS (VTO=0.4 KP=432E-6 GAMMA=0.2 PHI=.88)
.model EEPMOS PMOS (VTO=-0.4 KP=122E-6 GAMMA=0.2 PHI=.88)

.subckt myamp in_ out vdd vss

R0 vdd out 5000
MN0 out in_ vss vss EENMOS w=0.4u l=0.1u
C0 out vss 20n

.ends
