

/***********
* template made quickly by Daniel
* For demoing the rx with a slicer
***********/

// the declaratino comes straight from one of Byong's templates
module comparator1 #(
// parameters here
  
) (
  