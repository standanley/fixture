module my_inv (input in_, output out);
assign out = in_;
endmodule

