* Automatically generated file.
.include /home/dstanley/research/fixture/test_tsmc/phase_blender.spf
X0 ph_in[0] ph_in[1] ph_out thm_sel_bld[15] thm_sel_bld[14] thm_sel_bld[13] thm_sel_bld[12] thm_sel_bld[11] thm_sel_bld[10] thm_sel_bld[9] thm_sel_bld[8] thm_sel_bld[7] thm_sel_bld[6] thm_sel_bld[5] thm_sel_bld[4] thm_sel_bld[3] thm_sel_bld[2] thm_sel_bld[1] thm_sel_bld[0] phase_blender
.subckt inout_sw_mod sw_p sw_n ctl_p ctl_n
    G1 sw_p sw_n VCR PWL(1) ctl_p ctl_n 0v,1000000000.0 1v,1
.ends
X2 __ph_in[0]_v ph_in[0] __ph_in[0]_s 0 inout_sw_mod
V3 __ph_in[0]_v 0 DC 0 PWL(0 0 5.2001840282579426e-06 0 5.200384028257942e-06 0 5.500000000000001e-06 0 5.5002e-06 1 6.000000000000001e-06 1 6.000200000000001e-06 0 6.500000000000001e-06 0 6.500200000000001e-06 1 7.000000000000001e-06 1 7.0002e-06 0 7.500000000000001e-06 0 7.500200000000001e-06 1 8.000000000000001e-06 1 8.000200000000002e-06 0 8.500000000000002e-06 0 8.500200000000002e-06 1 9.000000000000002e-06 1 9.000200000000002e-06 0 9.500000000000004e-06 0 9.500200000000004e-06 1 1.0000000000000006e-05 1 1.0000200000000006e-05 0 1.0200184028257948e-05 0 1.0200384028257949e-05 0 1.540039991059075e-05 0 1.540059991059075e-05 0 1.570018402825795e-05 0 1.570038402825795e-05 1 1.6200184028257948e-05 1 1.620038402825795e-05 0 1.6700184028257947e-05 0 1.6700384028257947e-05 1 1.7200184028257945e-05 1 1.7200384028257946e-05 0 1.7700184028257944e-05 0 1.7700384028257944e-05 1 1.8200184028257943e-05 1 1.8200384028257943e-05 0 1.870018402825794e-05 0 1.870038402825794e-05 1 1.920018402825794e-05 1 1.920038402825794e-05 0 1.970018402825794e-05 0 1.970038402825794e-05 1 2.0200184028257937e-05 1 2.0200384028257937e-05 0 2.0400399910590735e-05 0 2.0400599910590735e-05 0 2.5600911580126338e-05 0 2.5601111580126338e-05 0 2.5900399910590733e-05 0 2.5900599910590733e-05 1 2.640039991059073e-05 1 2.6400599910590732e-05 0 2.690039991059073e-05 0 2.690059991059073e-05 1 2.740039991059073e-05 1 2.740059991059073e-05 0 2.7900399910590727e-05 0 2.7900599910590728e-05 1 2.8400399910590726e-05 1 2.8400599910590726e-05 0 2.8900399910590724e-05 0 2.8900599910590725e-05 1 2.9400399910590723e-05 1 2.9400599910590723e-05 0 2.990039991059072e-05 0 2.9900599910590722e-05 1 3.040039991059072e-05 1 3.040059991059072e-05 0 3.0600911580126324e-05 0 3.0601111580126324e-05 0 3.580158374751403e-05 0 3.580178374751403e-05 0 3.610091158012632e-05 0 3.610111158012632e-05 1 3.660091158012632e-05 1 3.660111158012632e-05 0 3.710091158012632e-05 0 3.710111158012632e-05 1 3.760091158012632e-05 1 3.760111158012632e-05 0 3.8100911580126316e-05 0 3.8101111580126317e-05 1 3.8600911580126315e-05 1 3.8601111580126315e-05 0 3.910091158012631e-05 0 3.9101111580126314e-05 1 3.960091158012631e-05 1 3.960111158012631e-05 0 4.010091158012631e-05 0 4.010111158012631e-05 1 4.060091158012631e-05 1 4.060111158012631e-05 0 4.080158374751402e-05 0 4.080178374751402e-05 0 4.60023907314374e-05 0 4.6002590731437404e-05 0 4.630158374751402e-05 0 4.630178374751402e-05 1 4.680158374751402e-05 1 4.680178374751402e-05 0 4.730158374751402e-05 0 4.730178374751402e-05 1 4.7801583747514016e-05 1 4.780178374751402e-05 0 4.8301583747514015e-05 0 4.8301783747514015e-05 1 4.8801583747514014e-05 1 4.8801783747514014e-05 0 4.930158374751401e-05 0 4.930178374751401e-05 1 4.980158374751401e-05 1 4.980178374751401e-05 0 5.030158374751401e-05 0 5.030178374751401e-05 1 5.080158374751401e-05 1 5.080178374751401e-05 0 5.10023907314374e-05 0 5.10025907314374e-05 0 5.6203456879677744e-05 0 5.6203656879677744e-05 0 5.65023907314374e-05 0 5.65025907314374e-05 1 5.70023907314374e-05 1 5.70025907314374e-05 0 5.75023907314374e-05 0 5.75025907314374e-05 1 5.80023907314374e-05 1 5.80025907314374e-05 0 5.8502390731437395e-05 0 5.8502590731437396e-05 1 5.9002390731437394e-05 1 5.9002590731437394e-05 0 5.950239073143739e-05 0 5.950259073143739e-05 1 6.000239073143739e-05 1 6.000259073143739e-05 0 6.050239073143739e-05 0 6.050259073143739e-05 1 6.100239073143739e-05 1 6.100259073143739e-05 0 6.120345687967774e-05 0 6.120365687967774e-05 0 6.640480297716098e-05 0 6.640500297716098e-05 0 6.670345687967774e-05 0 6.670365687967774e-05 1 6.720345687967773e-05 1 6.720365687967773e-05 0 6.770345687967771e-05 0 6.770365687967771e-05 1 6.82034568796777e-05 1 6.82036568796777e-05 0 6.870345687967768e-05 0 6.870365687967768e-05 1 6.920345687967767e-05 1 6.920365687967767e-05 0 6.970345687967765e-05 0 6.970365687967765e-05 1 7.020345687967764e-05 1 7.020365687967764e-05 0 7.070345687967762e-05 0 7.070365687967762e-05 1 7.120345687967761e-05 1 7.120365687967761e-05 0 7.140480297716086e-05 0 7.140500297716086e-05 0 7.660630340083568e-05 0 7.660650340083568e-05 0 7.690480297716086e-05 0 7.690500297716086e-05 1 7.740480297716086e-05 1 7.740500297716086e-05 0 7.790480297716086e-05 0 7.790500297716086e-05 1 7.840480297716085e-05 1 7.840500297716085e-05 0 7.890480297716085e-05 0 7.890500297716085e-05 1 7.940480297716085e-05 1 7.940500297716085e-05 0 7.990480297716085e-05 0 7.990500297716085e-05 1 8.040480297716085e-05 1 8.040500297716085e-05 0 8.090480297716085e-05 0 8.090500297716085e-05 1 8.140480297716085e-05 1 8.140500297716085e-05 0 8.160630340083568e-05 0 8.160650340083568e-05 0 8.68080003149639e-05 0 8.68082003149639e-05 0 8.71063034008357e-05 0 8.71065034008357e-05 1 8.760630340083568e-05 1 8.760650340083568e-05 0 8.810630340083566e-05 0 8.810650340083566e-05 1 8.860630340083565e-05 1 8.860650340083565e-05 0 8.910630340083563e-05 0 8.910650340083563e-05 1 8.960630340083562e-05 1 8.960650340083562e-05 0 9.01063034008356e-05 0 9.01065034008356e-05 1 9.060630340083559e-05 1 9.060650340083559e-05 0 9.110630340083557e-05 0 9.110650340083557e-05 1 9.160630340083556e-05 1 9.160650340083556e-05 0 9.180800031496378e-05 0 9.180820031496378e-05 0 9.700984556640298e-05 0 9.701004556640298e-05 0 9.730800031496379e-05 0 9.730820031496379e-05 1 9.78080003149638e-05 1 9.78082003149638e-05 0 9.830800031496382e-05 0 9.830820031496382e-05 1 9.880800031496383e-05 1 9.880820031496383e-05 0 9.930800031496384e-05 0 9.930820031496384e-05 1 9.980800031496385e-05 1 9.980820031496385e-05 0 0.00010030800031496386 0 0.00010030820031496386 1 0.00010080800031496388 1 0.00010080820031496388 0 0.00010130800031496389 0 0.00010130820031496389 1 0.0001018080003149639 1 0.0001018082003149639 0 0.00010200984556640312 0 0.00010201004556640312 0 0.00010721189158154771 0 0.00010721209158154771 0 0.00010750984556640313 0 0.00010751004556640313 1 0.00010800984556640311 1 0.00010801004556640311 0 0.0001085098455664031 0 0.0001085100455664031 1 0.00010900984556640308 1 0.00010901004556640308 0 0.00010950984556640307 0 0.00010951004556640307 1 0.00011000984556640305 1 0.00011001004556640305 0 0.00011050984556640304 0 0.00011051004556640304 1 0.00011100984556640302 1 0.00011101004556640302 0 0.00011150984556640301 0 0.00011151004556640301 1 0.00011200984556640299 1 0.00011201004556640299 0 0.00011221189158154759 0 0.00011221209158154759 0 0.00011741412374722472 0 0.00011741432374722472 0 0.00011771189158154758 0 0.00011771209158154758 1 0.00011821189158154756 1 0.00011821209158154756 0 0.00011871189158154755 0 0.00011871209158154755 1 0.00011921189158154753 1 0.00011921209158154753 0 0.00011971189158154752 0 0.00011971209158154752 1 0.0001202118915815475 1 0.0001202120915815475 0 0.00012071189158154749 0 0.00012071209158154749 1 0.00012121189158154747 1 0.00012121209158154747 0 0.00012171189158154747 0 0.00012171209158154747 1 0.00012221189158154747 1 0.00012221209158154746 0 0.0001224141237472246 0 0.00012241432374722458 0 0.00012761667966227716 0 0.00012761687966227715 0 0.00012791412374722462 0 0.0001279143237472246 1 0.00012841412374722463 1 0.00012841432374722462 0 0.00012891412374722465 0 0.00012891432374722463 1 0.00012941412374722466 1 0.00012941432374722464 0 0.00012991412374722467 0 0.00012991432374722466 1 0.00013041412374722468 1 0.00013041432374722467 0 0.0001309141237472247 0 0.00013091432374722468 1 0.0001314141237472247 1 0.0001314143237472247 0 0.00013191412374722472 0 0.0001319143237472247 1 0.00013241412374722473 1 0.00013241432374722472 0 0.0001326166796622773 0 0.0001326168796622773 0 0.00013781929267817238 0 0.00013781949267817236 0 0.00013811667966227734 0 0.00013811687966227732 1 0.00013861667966227735 1 0.00013861687966227733 0 0.00013911667966227736 0 0.00013911687966227735 1 0.00013961667966227737 1 0.00013961687966227736 0 0.00014011667966227738 0 0.00014011687966227737 1 0.0001406166796622774 1 0.00014061687966227738 0 0.0001411166796622774 0 0.0001411168796622774 1 0.00014161667966227742 1 0.0001416168796622774 0 0.00014211667966227743 0 0.00014211687966227742 1 0.00014261667966227745 1 0.00014261687966227743 0 0.00014281929267817253 0 0.0001428194926781725 0 0.000148022148519013 0 0.00014802234851901298 0 0.00014831929267817252 0 0.0001483194926781725 1 0.00014881929267817254 1 0.00014881949267817252 0 0.00014931929267817255 0 0.00014931949267817254 1 0.00014981929267817256 1 0.00014981949267817255 0 0.00015031929267817257 0 0.00015031949267817256 1 0.00015081929267817258 1 0.00015081949267817257 0 0.0001513192926781726 0 0.00015131949267817258 1 0.0001518192926781726 1 0.0001518194926781726 0 0.00015231929267817262 0 0.0001523194926781726 1 0.00015281929267817263 1 0.00015281949267817262 0 0.00015302214851901311 0 0.0001530223485190131 0 0.000158225310832565 0 0.00015822551083256498 0 0.0001585221485190131 0 0.0001585223485190131 1 0.00015902214851901312 1 0.0001590223485190131 0 0.00015952214851901314 0 0.00015952234851901312 1 0.00016002214851901315 1 0.00016002234851901314 0 0.00016052214851901316 0 0.00016052234851901315 1 0.00016102214851901317 1 0.00016102234851901316 0 0.00016152214851901319 0 0.00016152234851901317 1 0.0001620221485190132 1 0.00016202234851901318 0 0.0001625221485190132 0 0.0001625223485190132 1 0.00016302214851901322 1 0.0001630223485190132 0 0.00016322531083256511 0 0.0001632255108325651 0 0.0001684286310398012 0 0.0001684288310398012 0 0.00016872531083256514 0 0.00016872551083256513 1 0.00016922531083256512 1 0.0001692255108325651 0 0.00016972531083256514 0 0.00016972551083256512 1 0.00017022531083256515 1 0.00017022551083256514 0 0.00017072531083256516 0 0.00017072551083256515 1 0.00017122531083256517 1 0.00017122551083256516 0 0.00017172531083256519 0 0.00017172551083256517 1 0.0001722253108325652 1 0.00017222551083256518 0 0.0001727253108325652 0 0.0001727255108325652 1 0.00017322531083256522 1 0.0001732255108325652 0 0.0001734286310398013 0 0.00017342883103980129 0 0.00017863213915402182 0 0.0001786323391540218 0 0.00017892863103980132 0 0.0001789288310398013 1 0.00017942863103980134 1 0.00017942883103980132 0 0.00017992863103980135 0 0.00017992883103980134 1 0.00018042863103980136 1 0.00018042883103980135 0 0.00018092863103980137 0 0.00018092883103980136 1 0.00018142863103980138 1 0.00018142883103980137 0 0.0001819286310398014 0 0.00018192883103980138 1 0.0001824286310398014 1 0.0001824288310398014 0 0.00018292863103980142 0 0.0001829288310398014 1 0.00018342863103980143 1 0.00018342883103980142 0 0.00018363213915402194 0 0.00018363233915402193 0 0.0001888358186013159 0 0.0001888360186013159 0 0.00018913213915402197 0 0.00018913233915402196 1 0.00018963213915402198 1 0.00018963233915402197 0 0.000190132139154022 0 0.00019013233915402198 1 0.000190632139154022 1 0.000190632339154022 0 0.00019113213915402202 0 0.000191132339154022 1 0.00019163213915402203 1 0.00019163233915402202 0 0.00019213213915402204 0 0.00019213233915402203 1 0.00019263213915402205 1 0.00019263233915402204 0 0.00019313213915402207 0 0.00019313233915402205 1 0.00019363213915402208 1 0.00019363233915402206 0 0.00019383581860131602 0 0.000193836018601316 0 0.00019903971249211137 0 0.00019903991249211136 0 0.00019933581860131605 0 0.00019933601860131603 1 0.00019983581860131606 1 0.00019983601860131605 0 0.00020033581860131607 0 0.00020033601860131606 1 0.00020083581860131608 1 0.00020083601860131607 0 0.0002013358186013161 0 0.00020133601860131608 1 0.0002018358186013161 1 0.0002018360186013161 0 0.00020233581860131612 0 0.0002023360186013161 1 0.00020283581860131613 1 0.00020283601860131612 0 0.00020333581860131614 0 0.00020333601860131613 1 0.00020383581860131616 1 0.00020383601860131614 0 0.00020403971249211152 0 0.0002040399124921115 0 0.0002092437273079041 0 0.0002092439273079041 0 0.00020953971249211155 0 0.00020953991249211153 1 0.00021003971249211156 1 0.00021003991249211155 0 0.00021053971249211157 0 0.00021053991249211156 1 0.00021103971249211158 1 0.00021103991249211157 0 0.0002115397124921116 0 0.00021153991249211158 1 0.0002120397124921116 1 0.0002120399124921116 0 0.00021253971249211162 0 0.0002125399124921116 1 0.00021303971249211163 1 0.00021303991249211162 0 0.00021353971249211165 0 0.00021353991249211163 1 0.00021403971249211166 1 0.00021403991249211164 0 0.00021424372730790425 0 0.00021424392730790424 0 0.00021944808721675776 0 0.00021944828721675775 0 0.00021974372730790428 0 0.00021974392730790426 1 0.0002202437273079043 1 0.00022024392730790428 0 0.0002207437273079043 0 0.0002207439273079043 1 0.00022124372730790431 1 0.0002212439273079043 0 0.00022174372730790433 0 0.0002217439273079043 1 0.00022224372730790434 1 0.00022224392730790433 0 0.00022274372730790435 0 0.00022274392730790434 1 0.00022324372730790436 1 0.00022324392730790435 0 0.00022374372730790438 0 0.00022374392730790436 1 0.0002242437273079044 1 0.00022424392730790437 0 0.00022444808721675788 0 0.00022444828721675787 0 0.00022965261116331256 0 0.00022965281116331255 0 0.0002299480872167579 0 0.0002299482872167579 1 0.00023044808721675792 1 0.0002304482872167579 0 0.00023094808721675793 0 0.00023094828721675792 1 0.00023144808721675794 1 0.00023144828721675793 0 0.00023194808721675795 0 0.00023194828721675794 1 0.00023244808721675797 1 0.00023244828721675795 0 0.00023294808721675798 0 0.00023294828721675797 1 0.000233448087216758 1 0.00023344828721675798 0 0.000233948087216758 0 0.000233948287216758 1 0.00023444808721675802 1 0.000234448287216758 0 0.00023465261116331268 0 0.00023465281116331267 0 0.00023985725348777873 0 0.00023985745348777872 0 0.0002401526111633127 0 0.0002401528111633127 1 0.00024065261116331272 1 0.0002406528111633127 0 0.00024115261116331273 0 0.00024115281116331272 1 0.00024165261116331274 1 0.00024165281116331273 0 0.00024215261116331276 0 0.00024215281116331274 1 0.00024265261116331277 1 0.00024265281116331276 0 0.00024315261116331278 0 0.00024315281116331277 1 0.0002436526111633128 1 0.00024365281116331278 0 0.0002441526111633128 0 0.0002441528111633128 1 0.0002446526111633128 1 0.00024465281116331283 0 0.0002448572534877788 0 0.0002448574534877788 0 0.00025006213249421645 0 0.00025006233249421646 0 0.0002503572534877788 0 0.00025035745348777884 1 0.00025085725348777884 1 0.00025085745348777885 0 0.00025135725348777885 0 0.00025135745348777886 1 0.00025185725348777886 1 0.0002518574534877789 0 0.0002523572534877789 0 0.0002523574534877789 1 0.0002528572534877789 1 0.0002528574534877789 0 0.0002533572534877789 0 0.0002533574534877789 1 0.0002538572534877789 1 0.0002538574534877789 0 0.0002543572534877789 0 0.00025435745348777894 1 0.00025485725348777893 1 0.00025485745348777895 0 0.00025506213249421646 0 0.0002550623324942165 0 0.00026026732409400484 0 0.00026026752409400486 0 0.00026056213249421643 0 0.00026056233249421645 1 0.0002610621324942165 1 0.0002610623324942165 0 0.00026156213249421657 0 0.0002615623324942166 1 0.00026206213249421663 1 0.00026206233249421665 0 0.0002625621324942167 0 0.0002625623324942167 1 0.00026306213249421677 1 0.0002630623324942168 0 0.00026356213249421683 0 0.00026356233249421685 1 0.0002640621324942169 1 0.0002640623324942169 0 0.00026456213249421697 0 0.000264562332494217 1 0.00026506213249421703 1 0.00026506233249421705 0 0.00026526732409400534 0 0.00026526752409400536 0 0.00027047253727422333 0 0.00027047273727422334 0 0.0002707673240940054 0 0.00027076752409400544 1 0.0002712673240940054 1 0.0002712675240940054 0 0.00027176732409400534 0 0.00027176752409400535 1 0.0002722673240940053 1 0.0002722675240940053 0 0.00027276732409400525 0 0.00027276752409400527 1 0.0002732673240940052 1 0.0002732675240940052 0 0.00027376732409400517 0 0.0002737675240940052 1 0.00027426732409400513 1 0.00027426752409400514 0 0.0002747673240940051 0 0.0002747675240940051 1 0.00027526732409400504 1 0.00027526752409400506 0 0.00027547253727422285 0 0.00027547273727422287 0 0.0002806781009094726 0 0.0002806783009094726 0 0.0002809725372742229 0 0.0002809727372742229 1 0.0002814725372742229 1 0.0002814727372742229 0 0.0002819725372742229 0 0.0002819727372742229 1 0.0002824725372742229 1 0.00028247273727422293 0 0.00028297253727422293 0 0.00028297273727422294 1 0.00028347253727422294 1 0.00028347273727422295 0 0.00028397253727422295 0 0.00028397273727422297 1 0.00028447253727422296 1 0.000284472737274223 0 0.000284972537274223 0 0.000284972737274223 1 0.000285472537274223 1 0.000285472737274223 0 0.0002856781009094726 0 0.0002856783009094726 0 0.0002908838383549405 0 0.0002908840383549405 0 0.00029117810090947263 0 0.00029117830090947264 1 0.0002916781009094726 1 0.0002916783009094726 0 0.00029217810090947254 0 0.00029217830090947256 1 0.0002926781009094725 1 0.0002926783009094725 0 0.00029317810090947246 0 0.0002931783009094725 1 0.0002936781009094724 1 0.00029367830090947243 0 0.0002941781009094724 0 0.0002941783009094724 1 0.00029467810090947233 1 0.00029467830090947235 0 0.0002951781009094723 0 0.0002951783009094723 1 0.00029567810090947225 1 0.00029567830090947226 0 0.00029588383835494 0 0.00029588403835494 0 0.0003010896923277906 0 0.00030108989232779064 0 0.00030138383835493995 0 0.00030138403835493996 1 0.0003018838383549399 1 0.0003018840383549399 0 0.00030238383835493987 0 0.0003023840383549399 1 0.0003028838383549398 1 0.00030288403835493984 0 0.0003033838383549398 0 0.0003033840383549398 1 0.00030388383835493974 1 0.00030388403835493975 0 0.0003043838383549397 0 0.0003043840383549397 1 0.00030488383835493966 1 0.00030488403835493967 0 0.0003053838383549396 0 0.00030538403835493963 1 0.00030588383835493957 1 0.0003058840383549396 0 0.0003060896923277901 0 0.0003060898923277901 0 0.0003112957259554461 0 0.0003112959259554461 0 0.00031158969232779007 0 0.0003115898923277901 1 0.00031208969232779 1 0.00031208989232779004 0 0.00031258969232779 0 0.00031258989232779 1 0.00031308969232778994 1 0.00031308989232778996 0 0.0003135896923277899 0 0.0003135898923277899 1 0.00031408969232778986 1 0.00031408989232778987 0 0.0003145896923277898 0 0.00031458989232778983 1 0.0003150896923277898 1 0.0003150898923277898 0 0.00031558969232778973 0 0.00031558989232778975 1 0.0003160896923277897 1 0.0003160898923277897 0 0.00031629572595544557 0 0.0003162959259554456 0 0.0003215020377403174 0 0.00032150223774031744 0 0.00032179572595544554 0 0.00032179592595544556 1 0.0003222957259554456 1 0.0003222959259554456 0 0.0003227957259554457 0 0.0003227959259554457 1 0.00032329572595544574 1 0.00032329592595544576 0 0.0003237957259554458 0 0.0003237959259554458 1 0.0003242957259554459 1 0.0003242959259554459 0 0.00032479572595544594 0 0.00032479592595544595 1 0.000325295725955446 1 0.000325295925955446 0 0.0003257957259554461 0 0.0003257959259554461 1 0.00032629572595544614 1 0.00032629592595544615 0 0.0003265020377403179 0 0.00032650223774031794 0 0.0003317084673472993 0 0.00033170866734729933 0 0.000332002037740318 0 0.000332002237740318 1 0.00033250203774031807 1 0.0003325022377403181 0 0.00033300203774031813 0 0.00033300223774031815 1 0.0003335020377403182 1 0.0003335022377403182 0 0.00033400203774031827 0 0.0003340022377403183 1 0.00033450203774031833 1 0.00033450223774031835 0 0.0003350020377403184 0 0.0003350022377403184 1 0.00033550203774031847 1 0.0003355022377403185 0 0.00033600203774031853 0 0.00033600223774031855 1 0.0003365020377403186 1 0.0003365022377403186 0 0.00033670846734729987 0 0.0003367086673472999 0 0.000341915233652557 0 0.000341915433652557 0 0.00034220846734729984 0 0.00034220866734729986 1 0.0003427084673472998 1 0.0003427086673472998 0 0.00034320846734729976 0 0.0003432086673472998 1 0.0003437084673472997 1 0.00034370866734729973 0 0.0003442084673472997 0 0.0003442086673472997 1 0.00034470846734729963 1 0.00034470866734729965 0 0.0003452084673472996 0 0.0003452086673472996 1 0.00034570846734729955 1 0.00034570866734729956 0 0.0003462084673472995 0 0.0003462086673472995 1 0.00034670846734729947 1 0.0003467086673472995 0 0.00034691523365255644 0 0.00034691543365255646 0 0.00035212205306404026 0 0.0003521222530640403 0 0.0003524152336525565 0 0.00035241543365255654 1 0.0003529152336525565 1 0.0003529154336525565 0 0.00035341523365255644 0 0.00035341543365255645 1 0.0003539152336525564 1 0.0003539154336525564 0 0.00035441523365255636 0 0.00035441543365255637 1 0.0003549152336525563 1 0.00035491543365255633 0 0.00035541523365255627 0 0.0003554154336525563 1 0.00035591523365255623 1 0.00035591543365255624 0 0.0003564152336525562 0 0.0003564154336525562 1 0.00035691523365255615 1 0.00035691543365255616 0 0.0003571220530640398 0 0.0003571222530640398 0 0.00036232924646941806 0 0.00036232944646941807 0 0.0003626220530640398 0 0.00036262225306403983 1 0.0003631220530640398 1 0.00036312225306403984 0 0.00036362205306403984 0 0.00036362225306403985 1 0.00036412205306403985 1 0.00036412225306403986 0 0.00036462205306403986 0 0.0003646222530640399 1 0.0003651220530640399 1 0.0003651222530640399 0 0.0003656220530640399 0 0.0003656222530640399 1 0.0003661220530640399 1 0.0003661222530640399 0 0.0003666220530640399 0 0.0003666222530640399 1 0.0003671220530640399 1 0.00036712225306403994 0 0.00036732924646941807 0 0.0003673294464694181 0 0.0003725365334006625 0 0.0003725367334006625 0 0.0003728292464694181 0 0.0003728294464694181 1 0.0003733292464694181 1 0.0003733294464694181 0 0.0003738292464694181 0 0.00037382944646941813 1 0.00037432924646941813 1 0.00037432944646941814 0 0.00037482924646941814 0 0.00037482944646941816 1 0.00037532924646941816 1 0.00037532944646941817 0 0.00037582924646941817 0 0.0003758294464694182 1 0.0003763292464694182 1 0.0003763294464694182 0 0.0003768292464694182 0 0.0003768294464694182 1 0.0003773292464694182 1 0.0003773294464694182 0 0.0003775365334006625 0 0.0003775367334006625 0 0.00038274395561190434 0 0.00038274415561190435 0 0.0003830365334006625 0 0.00038303673340066253 1 0.0003835365334006625 1 0.0003835367334006625 0 0.00038403653340066243 0 0.00038403673340066245 1 0.0003845365334006624 1 0.0003845367334006624 0 0.00038503653340066235 0 0.00038503673340066236 1 0.0003855365334006623 1 0.0003855367334006623 0 0.00038603653340066226 0 0.0003860367334006623 1 0.0003865365334006622 1 0.00038653673340066224 0 0.0003870365334006622 0 0.0003870367334006622 1 0.00038753653340066214 1 0.00038753673340066215 0 0.0003877439556119038 0 0.0003877441556119038 0 0.00039295175422431375 0 0.00039295195422431377 0 0.00039324395561190383 0 0.00039324415561190385 1 0.00039374395561190384 1 0.00039374415561190386 0 0.00039424395561190386 0 0.00039424415561190387 1 0.00039474395561190387 1 0.0003947441556119039 0 0.0003952439556119039 0 0.0003952441556119039 1 0.0003957439556119039 1 0.0003957441556119039 0 0.0003962439556119039 0 0.0003962441556119039 1 0.0003967439556119039 1 0.00039674415561190393 0 0.00039724395561190393 0 0.00039724415561190394 1 0.00039774395561190394 1 0.00039774415561190396 0 0.00039795175422431377 0 0.0003979519542243138 0 0.00040315970887468036 0 0.00040315990887468037 0 0.00040345175422431385 0 0.00040345195422431386 1 0.0004039517542243139 1 0.0004039519542243139 0 0.000404451754224314 0 0.000404451954224314 1 0.00040495175422431405 1 0.00040495195422431406 0 0.0004054517542243141 0 0.0004054519542243141 1 0.0004059517542243142 1 0.0004059519542243142 0 0.00040645175422431424 0 0.00040645195422431426 1 0.0004069517542243143 1 0.0004069519542243143 0 0.0004074517542243144 0 0.0004074519542243144 1 0.00040795175422431444 1 0.00040795195422431446 0 0.0004081597088746809 0 0.0004081599088746809 0 0.0004133678210077549 0 0.0004133680210077549 0 0.0004136597088746809 0 0.0004136599088746809 1 0.00041415970887468095 1 0.00041415990887468096 0 0.000414659708874681 0 0.00041465990887468103 1 0.0004151597088746811 1 0.0004151599088746811 0 0.00041565970887468115 0 0.00041565990887468116 1 0.0004161597088746812 1 0.00041615990887468123 0 0.0004166597088746813 0 0.0004166599088746813 1 0.00041715970887468135 1 0.00041715990887468136 0 0.0004176597088746814 0 0.00041765990887468143 1 0.0004181597088746815 1 0.0004181599088746815 0 0.0004183678210077554 0 0.0004183680210077554 0 0.00042357605238244213 0 0.00042357625238244215 0 0.0004238678210077554 0 0.0004238680210077554 1 0.0004243678210077554 1 0.00042436802100775543 0 0.00042486782100775543 0 0.00042486802100775544 1 0.00042536782100775544 1 0.00042536802100775546 0 0.00042586782100775545 0 0.00042586802100775547 1 0.00042636782100775547 1 0.0004263680210077555 0 0.0004268678210077555 0 0.0004268680210077555 1 0.0004273678210077555 1 0.0004273680210077555 0 0.0004278678210077555 0 0.0004278680210077555 1 0.0004283678210077555 1 0.00042836802100775553 0 0.00042857605238244215 0 0.00042857625238244216 0 0.0004337845821168645 0 0.00043378478211686454 0 0.00043407605238244217 0 0.0004340762523824422 1 0.00043457605238244224 1 0.00043457625238244225 0 0.0004350760523824423 0 0.0004350762523824423 1 0.00043557605238244237 1 0.0004355762523824424 0 0.00043607605238244244 0 0.00043607625238244245 1 0.0004365760523824425 1 0.0004365762523824425 0 0.00043707605238244257 0 0.0004370762523824426 1 0.00043757605238244263 1 0.00043757625238244265 0 0.0004380760523824427 0 0.0004380762523824427 1 0.00043857605238244277 1 0.0004385762523824428 0 0.000438784582116865 0 0.00043878478211686504 0 0.00044399329473837737 0 0.0004439934947383774 0 0.00044428458211686505 0 0.00044428478211686506 1 0.00044478458211686506 1 0.0004447847821168651 0 0.0004452845821168651 0 0.0004452847821168651 1 0.0004457845821168651 1 0.0004457847821168651 0 0.0004462845821168651 0 0.0004462847821168651 1 0.0004467845821168651 1 0.0004467847821168651 0 0.0004472845821168651 0 0.00044728478211686514 1 0.00044778458211686514 1 0.00044778478211686515 0 0.00044828458211686515 0 0.00044828478211686516 1 0.00044878458211686516 1 0.0004487847821168652 0 0.0004489932947383774 0 0.0004489934947383774 0 0.0004542021916109949 0 0.0004542023916109949 0 0.0004544932947383774 0 0.0004544934947383774 1 0.00045499329473837737 1 0.0004549934947383774 0 0.0004554932947383773 0 0.00045549349473837734 1 0.0004559932947383773 1 0.0004559934947383773 0 0.00045649329473837724 0 0.00045649349473837725 1 0.0004569932947383772 1 0.0004569934947383772 0 0.00045749329473837716 0 0.00045749349473837717 1 0.0004579932947383771 1 0.00045799349473837713 0 0.00045849329473837707 0 0.0004584934947383771 1 0.00045899329473837703 1 0.00045899349473837704 0 0.00045920219161099435 0 0.00045920239161099436 0 0.00046441127816508496 0 0.00046441147816508497 0 0.0004647021916109944 0 0.0004647023916109944 1 0.0004652021916109944 1 0.0004652023916109944 0 0.0004657021916109944 0 0.0004657023916109944 1 0.0004662021916109944 1 0.0004662023916109944 0 0.0004667021916109944 0 0.00046670239161099444 1 0.00046720219161099444 1 0.00046720239161099445 0 0.00046770219161099445 0 0.00046770239161099446 1 0.00046820219161099446 1 0.0004682023916109945 0 0.00046870219161099447 0 0.0004687023916109945 1 0.0004692021916109945 1 0.0004692023916109945 0 0.00046941127816508497 0 0.000469411478165085 0 0.0004746205704165872 0 0.0004746207704165872 0 0.000474911278165085 0 0.000474911478165085 1 0.00047541127816508506 1 0.0004754114781650851 0 0.0004759112781650851 0 0.00047591147816508514 1 0.0004764112781650852 1 0.0004764114781650852 0 0.00047691127816508526 0 0.0004769114781650853 1 0.0004774112781650853 1 0.00047741147816508534 0 0.0004779112781650854 0 0.0004779114781650854 1 0.00047841127816508546 1 0.00047841147816508547 0 0.0004789112781650855 0 0.00047891147816508554 1 0.00047941127816508554 1 0.00047941147816508555 0 0.00047962057041658765 0 0.00047962077041658767 0 0.00048483012515769053 0 0.00048483032515769055 0 0.0004851205704165877 0 0.0004851207704165877 1 0.0004856205704165877 1 0.0004856207704165877 0 0.0004861205704165877 0 0.0004861207704165877 1 0.0004866205704165877 1 0.00048662077041658773 0 0.00048712057041658773 0 0.00048712077041658774 1 0.00048762057041658774 1 0.00048762077041658775 0 0.00048812057041658775 0 0.00048812077041658777 1 0.0004886205704165877 1 0.0004886207704165877 0 0.0004891205704165878 0 0.0004891207704165877 1 0.0004896205704165878 1 0.0004896207704165878 0 0.0004898301251576905 0 0.0004898303251576905 0 0.000495039780822236 0 0.000495039980822236 0 0.0004953301251576906 0 0.0004953303251576906 1 0.0004958301251576906 1 0.0004958303251576905 0 0.0004963301251576906 0 0.0004963303251576906 1 0.0004968301251576907 1 0.0004968303251576907 0 0.0004973301251576908 0 0.0004973303251576907 1 0.0004978301251576908 1 0.0004978303251576908 0 0.0004983301251576909 0 0.0004983303251576909 1 0.000498830125157691 1 0.0004988303251576909 0 0.000499330125157691 0 0.000499330325157691 1 0.0004998301251576911 1 0.0004998303251576911 0 0.0005000397808222364 0 0.0005000399808222363 0 0.0005052496159810823 0 0.0005052498159810822 0 0.0005055397808222363 0 0.0005055399808222363 1 0.0005060397808222364 1 0.0005060399808222364 0 0.0005065397808222365 0 0.0005065399808222364 1 0.0005070397808222365 1 0.0005070399808222365 0 0.0005075397808222366 0 0.0005075399808222366 1 0.0005080397808222367 1 0.0005080399808222366 0 0.0005085397808222367 0 0.0005085399808222367 1 0.0005090397808222368 1 0.0005090399808222368 0 0.0005095397808222369 0 0.0005095399808222368 1 0.000510039780822237 1 0.0005100399808222369 0 0.0005102496159810827 0)
V4 __ph_in[0]_s 0 DC 1 PWL(0 1 5.2001840282579426e-06 1 5.200384028257942e-06 1 5.500000000000001e-06 1 5.5002e-06 1 6.000000000000001e-06 1 6.000200000000001e-06 1 6.500000000000001e-06 1 6.500200000000001e-06 1 7.000000000000001e-06 1 7.0002e-06 1 7.500000000000001e-06 1 7.500200000000001e-06 1 8.000000000000001e-06 1 8.000200000000002e-06 1 8.500000000000002e-06 1 8.500200000000002e-06 1 9.000000000000002e-06 1 9.000200000000002e-06 1 9.500000000000004e-06 1 9.500200000000004e-06 1 1.0000000000000006e-05 1 1.0000200000000006e-05 1 1.0200184028257948e-05 1 1.0200384028257949e-05 1 1.540039991059075e-05 1 1.540059991059075e-05 1 1.570018402825795e-05 1 1.570038402825795e-05 1 1.6200184028257948e-05 1 1.620038402825795e-05 1 1.6700184028257947e-05 1 1.6700384028257947e-05 1 1.7200184028257945e-05 1 1.7200384028257946e-05 1 1.7700184028257944e-05 1 1.7700384028257944e-05 1 1.8200184028257943e-05 1 1.8200384028257943e-05 1 1.870018402825794e-05 1 1.870038402825794e-05 1 1.920018402825794e-05 1 1.920038402825794e-05 1 1.970018402825794e-05 1 1.970038402825794e-05 1 2.0200184028257937e-05 1 2.0200384028257937e-05 1 2.0400399910590735e-05 1 2.0400599910590735e-05 1 2.5600911580126338e-05 1 2.5601111580126338e-05 1 2.5900399910590733e-05 1 2.5900599910590733e-05 1 2.640039991059073e-05 1 2.6400599910590732e-05 1 2.690039991059073e-05 1 2.690059991059073e-05 1 2.740039991059073e-05 1 2.740059991059073e-05 1 2.7900399910590727e-05 1 2.7900599910590728e-05 1 2.8400399910590726e-05 1 2.8400599910590726e-05 1 2.8900399910590724e-05 1 2.8900599910590725e-05 1 2.9400399910590723e-05 1 2.9400599910590723e-05 1 2.990039991059072e-05 1 2.9900599910590722e-05 1 3.040039991059072e-05 1 3.040059991059072e-05 1 3.0600911580126324e-05 1 3.0601111580126324e-05 1 3.580158374751403e-05 1 3.580178374751403e-05 1 3.610091158012632e-05 1 3.610111158012632e-05 1 3.660091158012632e-05 1 3.660111158012632e-05 1 3.710091158012632e-05 1 3.710111158012632e-05 1 3.760091158012632e-05 1 3.760111158012632e-05 1 3.8100911580126316e-05 1 3.8101111580126317e-05 1 3.8600911580126315e-05 1 3.8601111580126315e-05 1 3.910091158012631e-05 1 3.9101111580126314e-05 1 3.960091158012631e-05 1 3.960111158012631e-05 1 4.010091158012631e-05 1 4.010111158012631e-05 1 4.060091158012631e-05 1 4.060111158012631e-05 1 4.080158374751402e-05 1 4.080178374751402e-05 1 4.60023907314374e-05 1 4.6002590731437404e-05 1 4.630158374751402e-05 1 4.630178374751402e-05 1 4.680158374751402e-05 1 4.680178374751402e-05 1 4.730158374751402e-05 1 4.730178374751402e-05 1 4.7801583747514016e-05 1 4.780178374751402e-05 1 4.8301583747514015e-05 1 4.8301783747514015e-05 1 4.8801583747514014e-05 1 4.8801783747514014e-05 1 4.930158374751401e-05 1 4.930178374751401e-05 1 4.980158374751401e-05 1 4.980178374751401e-05 1 5.030158374751401e-05 1 5.030178374751401e-05 1 5.080158374751401e-05 1 5.080178374751401e-05 1 5.10023907314374e-05 1 5.10025907314374e-05 1 5.6203456879677744e-05 1 5.6203656879677744e-05 1 5.65023907314374e-05 1 5.65025907314374e-05 1 5.70023907314374e-05 1 5.70025907314374e-05 1 5.75023907314374e-05 1 5.75025907314374e-05 1 5.80023907314374e-05 1 5.80025907314374e-05 1 5.8502390731437395e-05 1 5.8502590731437396e-05 1 5.9002390731437394e-05 1 5.9002590731437394e-05 1 5.950239073143739e-05 1 5.950259073143739e-05 1 6.000239073143739e-05 1 6.000259073143739e-05 1 6.050239073143739e-05 1 6.050259073143739e-05 1 6.100239073143739e-05 1 6.100259073143739e-05 1 6.120345687967774e-05 1 6.120365687967774e-05 1 6.640480297716098e-05 1 6.640500297716098e-05 1 6.670345687967774e-05 1 6.670365687967774e-05 1 6.720345687967773e-05 1 6.720365687967773e-05 1 6.770345687967771e-05 1 6.770365687967771e-05 1 6.82034568796777e-05 1 6.82036568796777e-05 1 6.870345687967768e-05 1 6.870365687967768e-05 1 6.920345687967767e-05 1 6.920365687967767e-05 1 6.970345687967765e-05 1 6.970365687967765e-05 1 7.020345687967764e-05 1 7.020365687967764e-05 1 7.070345687967762e-05 1 7.070365687967762e-05 1 7.120345687967761e-05 1 7.120365687967761e-05 1 7.140480297716086e-05 1 7.140500297716086e-05 1 7.660630340083568e-05 1 7.660650340083568e-05 1 7.690480297716086e-05 1 7.690500297716086e-05 1 7.740480297716086e-05 1 7.740500297716086e-05 1 7.790480297716086e-05 1 7.790500297716086e-05 1 7.840480297716085e-05 1 7.840500297716085e-05 1 7.890480297716085e-05 1 7.890500297716085e-05 1 7.940480297716085e-05 1 7.940500297716085e-05 1 7.990480297716085e-05 1 7.990500297716085e-05 1 8.040480297716085e-05 1 8.040500297716085e-05 1 8.090480297716085e-05 1 8.090500297716085e-05 1 8.140480297716085e-05 1 8.140500297716085e-05 1 8.160630340083568e-05 1 8.160650340083568e-05 1 8.68080003149639e-05 1 8.68082003149639e-05 1 8.71063034008357e-05 1 8.71065034008357e-05 1 8.760630340083568e-05 1 8.760650340083568e-05 1 8.810630340083566e-05 1 8.810650340083566e-05 1 8.860630340083565e-05 1 8.860650340083565e-05 1 8.910630340083563e-05 1 8.910650340083563e-05 1 8.960630340083562e-05 1 8.960650340083562e-05 1 9.01063034008356e-05 1 9.01065034008356e-05 1 9.060630340083559e-05 1 9.060650340083559e-05 1 9.110630340083557e-05 1 9.110650340083557e-05 1 9.160630340083556e-05 1 9.160650340083556e-05 1 9.180800031496378e-05 1 9.180820031496378e-05 1 9.700984556640298e-05 1 9.701004556640298e-05 1 9.730800031496379e-05 1 9.730820031496379e-05 1 9.78080003149638e-05 1 9.78082003149638e-05 1 9.830800031496382e-05 1 9.830820031496382e-05 1 9.880800031496383e-05 1 9.880820031496383e-05 1 9.930800031496384e-05 1 9.930820031496384e-05 1 9.980800031496385e-05 1 9.980820031496385e-05 1 0.00010030800031496386 1 0.00010030820031496386 1 0.00010080800031496388 1 0.00010080820031496388 1 0.00010130800031496389 1 0.00010130820031496389 1 0.0001018080003149639 1 0.0001018082003149639 1 0.00010200984556640312 1 0.00010201004556640312 1 0.00010721189158154771 1 0.00010721209158154771 1 0.00010750984556640313 1 0.00010751004556640313 1 0.00010800984556640311 1 0.00010801004556640311 1 0.0001085098455664031 1 0.0001085100455664031 1 0.00010900984556640308 1 0.00010901004556640308 1 0.00010950984556640307 1 0.00010951004556640307 1 0.00011000984556640305 1 0.00011001004556640305 1 0.00011050984556640304 1 0.00011051004556640304 1 0.00011100984556640302 1 0.00011101004556640302 1 0.00011150984556640301 1 0.00011151004556640301 1 0.00011200984556640299 1 0.00011201004556640299 1 0.00011221189158154759 1 0.00011221209158154759 1 0.00011741412374722472 1 0.00011741432374722472 1 0.00011771189158154758 1 0.00011771209158154758 1 0.00011821189158154756 1 0.00011821209158154756 1 0.00011871189158154755 1 0.00011871209158154755 1 0.00011921189158154753 1 0.00011921209158154753 1 0.00011971189158154752 1 0.00011971209158154752 1 0.0001202118915815475 1 0.0001202120915815475 1 0.00012071189158154749 1 0.00012071209158154749 1 0.00012121189158154747 1 0.00012121209158154747 1 0.00012171189158154747 1 0.00012171209158154747 1 0.00012221189158154747 1 0.00012221209158154746 1 0.0001224141237472246 1 0.00012241432374722458 1 0.00012761667966227716 1 0.00012761687966227715 1 0.00012791412374722462 1 0.0001279143237472246 1 0.00012841412374722463 1 0.00012841432374722462 1 0.00012891412374722465 1 0.00012891432374722463 1 0.00012941412374722466 1 0.00012941432374722464 1 0.00012991412374722467 1 0.00012991432374722466 1 0.00013041412374722468 1 0.00013041432374722467 1 0.0001309141237472247 1 0.00013091432374722468 1 0.0001314141237472247 1 0.0001314143237472247 1 0.00013191412374722472 1 0.0001319143237472247 1 0.00013241412374722473 1 0.00013241432374722472 1 0.0001326166796622773 1 0.0001326168796622773 1 0.00013781929267817238 1 0.00013781949267817236 1 0.00013811667966227734 1 0.00013811687966227732 1 0.00013861667966227735 1 0.00013861687966227733 1 0.00013911667966227736 1 0.00013911687966227735 1 0.00013961667966227737 1 0.00013961687966227736 1 0.00014011667966227738 1 0.00014011687966227737 1 0.0001406166796622774 1 0.00014061687966227738 1 0.0001411166796622774 1 0.0001411168796622774 1 0.00014161667966227742 1 0.0001416168796622774 1 0.00014211667966227743 1 0.00014211687966227742 1 0.00014261667966227745 1 0.00014261687966227743 1 0.00014281929267817253 1 0.0001428194926781725 1 0.000148022148519013 1 0.00014802234851901298 1 0.00014831929267817252 1 0.0001483194926781725 1 0.00014881929267817254 1 0.00014881949267817252 1 0.00014931929267817255 1 0.00014931949267817254 1 0.00014981929267817256 1 0.00014981949267817255 1 0.00015031929267817257 1 0.00015031949267817256 1 0.00015081929267817258 1 0.00015081949267817257 1 0.0001513192926781726 1 0.00015131949267817258 1 0.0001518192926781726 1 0.0001518194926781726 1 0.00015231929267817262 1 0.0001523194926781726 1 0.00015281929267817263 1 0.00015281949267817262 1 0.00015302214851901311 1 0.0001530223485190131 1 0.000158225310832565 1 0.00015822551083256498 1 0.0001585221485190131 1 0.0001585223485190131 1 0.00015902214851901312 1 0.0001590223485190131 1 0.00015952214851901314 1 0.00015952234851901312 1 0.00016002214851901315 1 0.00016002234851901314 1 0.00016052214851901316 1 0.00016052234851901315 1 0.00016102214851901317 1 0.00016102234851901316 1 0.00016152214851901319 1 0.00016152234851901317 1 0.0001620221485190132 1 0.00016202234851901318 1 0.0001625221485190132 1 0.0001625223485190132 1 0.00016302214851901322 1 0.0001630223485190132 1 0.00016322531083256511 1 0.0001632255108325651 1 0.0001684286310398012 1 0.0001684288310398012 1 0.00016872531083256514 1 0.00016872551083256513 1 0.00016922531083256512 1 0.0001692255108325651 1 0.00016972531083256514 1 0.00016972551083256512 1 0.00017022531083256515 1 0.00017022551083256514 1 0.00017072531083256516 1 0.00017072551083256515 1 0.00017122531083256517 1 0.00017122551083256516 1 0.00017172531083256519 1 0.00017172551083256517 1 0.0001722253108325652 1 0.00017222551083256518 1 0.0001727253108325652 1 0.0001727255108325652 1 0.00017322531083256522 1 0.0001732255108325652 1 0.0001734286310398013 1 0.00017342883103980129 1 0.00017863213915402182 1 0.0001786323391540218 1 0.00017892863103980132 1 0.0001789288310398013 1 0.00017942863103980134 1 0.00017942883103980132 1 0.00017992863103980135 1 0.00017992883103980134 1 0.00018042863103980136 1 0.00018042883103980135 1 0.00018092863103980137 1 0.00018092883103980136 1 0.00018142863103980138 1 0.00018142883103980137 1 0.0001819286310398014 1 0.00018192883103980138 1 0.0001824286310398014 1 0.0001824288310398014 1 0.00018292863103980142 1 0.0001829288310398014 1 0.00018342863103980143 1 0.00018342883103980142 1 0.00018363213915402194 1 0.00018363233915402193 1 0.0001888358186013159 1 0.0001888360186013159 1 0.00018913213915402197 1 0.00018913233915402196 1 0.00018963213915402198 1 0.00018963233915402197 1 0.000190132139154022 1 0.00019013233915402198 1 0.000190632139154022 1 0.000190632339154022 1 0.00019113213915402202 1 0.000191132339154022 1 0.00019163213915402203 1 0.00019163233915402202 1 0.00019213213915402204 1 0.00019213233915402203 1 0.00019263213915402205 1 0.00019263233915402204 1 0.00019313213915402207 1 0.00019313233915402205 1 0.00019363213915402208 1 0.00019363233915402206 1 0.00019383581860131602 1 0.000193836018601316 1 0.00019903971249211137 1 0.00019903991249211136 1 0.00019933581860131605 1 0.00019933601860131603 1 0.00019983581860131606 1 0.00019983601860131605 1 0.00020033581860131607 1 0.00020033601860131606 1 0.00020083581860131608 1 0.00020083601860131607 1 0.0002013358186013161 1 0.00020133601860131608 1 0.0002018358186013161 1 0.0002018360186013161 1 0.00020233581860131612 1 0.0002023360186013161 1 0.00020283581860131613 1 0.00020283601860131612 1 0.00020333581860131614 1 0.00020333601860131613 1 0.00020383581860131616 1 0.00020383601860131614 1 0.00020403971249211152 1 0.0002040399124921115 1 0.0002092437273079041 1 0.0002092439273079041 1 0.00020953971249211155 1 0.00020953991249211153 1 0.00021003971249211156 1 0.00021003991249211155 1 0.00021053971249211157 1 0.00021053991249211156 1 0.00021103971249211158 1 0.00021103991249211157 1 0.0002115397124921116 1 0.00021153991249211158 1 0.0002120397124921116 1 0.0002120399124921116 1 0.00021253971249211162 1 0.0002125399124921116 1 0.00021303971249211163 1 0.00021303991249211162 1 0.00021353971249211165 1 0.00021353991249211163 1 0.00021403971249211166 1 0.00021403991249211164 1 0.00021424372730790425 1 0.00021424392730790424 1 0.00021944808721675776 1 0.00021944828721675775 1 0.00021974372730790428 1 0.00021974392730790426 1 0.0002202437273079043 1 0.00022024392730790428 1 0.0002207437273079043 1 0.0002207439273079043 1 0.00022124372730790431 1 0.0002212439273079043 1 0.00022174372730790433 1 0.0002217439273079043 1 0.00022224372730790434 1 0.00022224392730790433 1 0.00022274372730790435 1 0.00022274392730790434 1 0.00022324372730790436 1 0.00022324392730790435 1 0.00022374372730790438 1 0.00022374392730790436 1 0.0002242437273079044 1 0.00022424392730790437 1 0.00022444808721675788 1 0.00022444828721675787 1 0.00022965261116331256 1 0.00022965281116331255 1 0.0002299480872167579 1 0.0002299482872167579 1 0.00023044808721675792 1 0.0002304482872167579 1 0.00023094808721675793 1 0.00023094828721675792 1 0.00023144808721675794 1 0.00023144828721675793 1 0.00023194808721675795 1 0.00023194828721675794 1 0.00023244808721675797 1 0.00023244828721675795 1 0.00023294808721675798 1 0.00023294828721675797 1 0.000233448087216758 1 0.00023344828721675798 1 0.000233948087216758 1 0.000233948287216758 1 0.00023444808721675802 1 0.000234448287216758 1 0.00023465261116331268 1 0.00023465281116331267 1 0.00023985725348777873 1 0.00023985745348777872 1 0.0002401526111633127 1 0.0002401528111633127 1 0.00024065261116331272 1 0.0002406528111633127 1 0.00024115261116331273 1 0.00024115281116331272 1 0.00024165261116331274 1 0.00024165281116331273 1 0.00024215261116331276 1 0.00024215281116331274 1 0.00024265261116331277 1 0.00024265281116331276 1 0.00024315261116331278 1 0.00024315281116331277 1 0.0002436526111633128 1 0.00024365281116331278 1 0.0002441526111633128 1 0.0002441528111633128 1 0.0002446526111633128 1 0.00024465281116331283 1 0.0002448572534877788 1 0.0002448574534877788 1 0.00025006213249421645 1 0.00025006233249421646 1 0.0002503572534877788 1 0.00025035745348777884 1 0.00025085725348777884 1 0.00025085745348777885 1 0.00025135725348777885 1 0.00025135745348777886 1 0.00025185725348777886 1 0.0002518574534877789 1 0.0002523572534877789 1 0.0002523574534877789 1 0.0002528572534877789 1 0.0002528574534877789 1 0.0002533572534877789 1 0.0002533574534877789 1 0.0002538572534877789 1 0.0002538574534877789 1 0.0002543572534877789 1 0.00025435745348777894 1 0.00025485725348777893 1 0.00025485745348777895 1 0.00025506213249421646 1 0.0002550623324942165 1 0.00026026732409400484 1 0.00026026752409400486 1 0.00026056213249421643 1 0.00026056233249421645 1 0.0002610621324942165 1 0.0002610623324942165 1 0.00026156213249421657 1 0.0002615623324942166 1 0.00026206213249421663 1 0.00026206233249421665 1 0.0002625621324942167 1 0.0002625623324942167 1 0.00026306213249421677 1 0.0002630623324942168 1 0.00026356213249421683 1 0.00026356233249421685 1 0.0002640621324942169 1 0.0002640623324942169 1 0.00026456213249421697 1 0.000264562332494217 1 0.00026506213249421703 1 0.00026506233249421705 1 0.00026526732409400534 1 0.00026526752409400536 1 0.00027047253727422333 1 0.00027047273727422334 1 0.0002707673240940054 1 0.00027076752409400544 1 0.0002712673240940054 1 0.0002712675240940054 1 0.00027176732409400534 1 0.00027176752409400535 1 0.0002722673240940053 1 0.0002722675240940053 1 0.00027276732409400525 1 0.00027276752409400527 1 0.0002732673240940052 1 0.0002732675240940052 1 0.00027376732409400517 1 0.0002737675240940052 1 0.00027426732409400513 1 0.00027426752409400514 1 0.0002747673240940051 1 0.0002747675240940051 1 0.00027526732409400504 1 0.00027526752409400506 1 0.00027547253727422285 1 0.00027547273727422287 1 0.0002806781009094726 1 0.0002806783009094726 1 0.0002809725372742229 1 0.0002809727372742229 1 0.0002814725372742229 1 0.0002814727372742229 1 0.0002819725372742229 1 0.0002819727372742229 1 0.0002824725372742229 1 0.00028247273727422293 1 0.00028297253727422293 1 0.00028297273727422294 1 0.00028347253727422294 1 0.00028347273727422295 1 0.00028397253727422295 1 0.00028397273727422297 1 0.00028447253727422296 1 0.000284472737274223 1 0.000284972537274223 1 0.000284972737274223 1 0.000285472537274223 1 0.000285472737274223 1 0.0002856781009094726 1 0.0002856783009094726 1 0.0002908838383549405 1 0.0002908840383549405 1 0.00029117810090947263 1 0.00029117830090947264 1 0.0002916781009094726 1 0.0002916783009094726 1 0.00029217810090947254 1 0.00029217830090947256 1 0.0002926781009094725 1 0.0002926783009094725 1 0.00029317810090947246 1 0.0002931783009094725 1 0.0002936781009094724 1 0.00029367830090947243 1 0.0002941781009094724 1 0.0002941783009094724 1 0.00029467810090947233 1 0.00029467830090947235 1 0.0002951781009094723 1 0.0002951783009094723 1 0.00029567810090947225 1 0.00029567830090947226 1 0.00029588383835494 1 0.00029588403835494 1 0.0003010896923277906 1 0.00030108989232779064 1 0.00030138383835493995 1 0.00030138403835493996 1 0.0003018838383549399 1 0.0003018840383549399 1 0.00030238383835493987 1 0.0003023840383549399 1 0.0003028838383549398 1 0.00030288403835493984 1 0.0003033838383549398 1 0.0003033840383549398 1 0.00030388383835493974 1 0.00030388403835493975 1 0.0003043838383549397 1 0.0003043840383549397 1 0.00030488383835493966 1 0.00030488403835493967 1 0.0003053838383549396 1 0.00030538403835493963 1 0.00030588383835493957 1 0.0003058840383549396 1 0.0003060896923277901 1 0.0003060898923277901 1 0.0003112957259554461 1 0.0003112959259554461 1 0.00031158969232779007 1 0.0003115898923277901 1 0.00031208969232779 1 0.00031208989232779004 1 0.00031258969232779 1 0.00031258989232779 1 0.00031308969232778994 1 0.00031308989232778996 1 0.0003135896923277899 1 0.0003135898923277899 1 0.00031408969232778986 1 0.00031408989232778987 1 0.0003145896923277898 1 0.00031458989232778983 1 0.0003150896923277898 1 0.0003150898923277898 1 0.00031558969232778973 1 0.00031558989232778975 1 0.0003160896923277897 1 0.0003160898923277897 1 0.00031629572595544557 1 0.0003162959259554456 1 0.0003215020377403174 1 0.00032150223774031744 1 0.00032179572595544554 1 0.00032179592595544556 1 0.0003222957259554456 1 0.0003222959259554456 1 0.0003227957259554457 1 0.0003227959259554457 1 0.00032329572595544574 1 0.00032329592595544576 1 0.0003237957259554458 1 0.0003237959259554458 1 0.0003242957259554459 1 0.0003242959259554459 1 0.00032479572595544594 1 0.00032479592595544595 1 0.000325295725955446 1 0.000325295925955446 1 0.0003257957259554461 1 0.0003257959259554461 1 0.00032629572595544614 1 0.00032629592595544615 1 0.0003265020377403179 1 0.00032650223774031794 1 0.0003317084673472993 1 0.00033170866734729933 1 0.000332002037740318 1 0.000332002237740318 1 0.00033250203774031807 1 0.0003325022377403181 1 0.00033300203774031813 1 0.00033300223774031815 1 0.0003335020377403182 1 0.0003335022377403182 1 0.00033400203774031827 1 0.0003340022377403183 1 0.00033450203774031833 1 0.00033450223774031835 1 0.0003350020377403184 1 0.0003350022377403184 1 0.00033550203774031847 1 0.0003355022377403185 1 0.00033600203774031853 1 0.00033600223774031855 1 0.0003365020377403186 1 0.0003365022377403186 1 0.00033670846734729987 1 0.0003367086673472999 1 0.000341915233652557 1 0.000341915433652557 1 0.00034220846734729984 1 0.00034220866734729986 1 0.0003427084673472998 1 0.0003427086673472998 1 0.00034320846734729976 1 0.0003432086673472998 1 0.0003437084673472997 1 0.00034370866734729973 1 0.0003442084673472997 1 0.0003442086673472997 1 0.00034470846734729963 1 0.00034470866734729965 1 0.0003452084673472996 1 0.0003452086673472996 1 0.00034570846734729955 1 0.00034570866734729956 1 0.0003462084673472995 1 0.0003462086673472995 1 0.00034670846734729947 1 0.0003467086673472995 1 0.00034691523365255644 1 0.00034691543365255646 1 0.00035212205306404026 1 0.0003521222530640403 1 0.0003524152336525565 1 0.00035241543365255654 1 0.0003529152336525565 1 0.0003529154336525565 1 0.00035341523365255644 1 0.00035341543365255645 1 0.0003539152336525564 1 0.0003539154336525564 1 0.00035441523365255636 1 0.00035441543365255637 1 0.0003549152336525563 1 0.00035491543365255633 1 0.00035541523365255627 1 0.0003554154336525563 1 0.00035591523365255623 1 0.00035591543365255624 1 0.0003564152336525562 1 0.0003564154336525562 1 0.00035691523365255615 1 0.00035691543365255616 1 0.0003571220530640398 1 0.0003571222530640398 1 0.00036232924646941806 1 0.00036232944646941807 1 0.0003626220530640398 1 0.00036262225306403983 1 0.0003631220530640398 1 0.00036312225306403984 1 0.00036362205306403984 1 0.00036362225306403985 1 0.00036412205306403985 1 0.00036412225306403986 1 0.00036462205306403986 1 0.0003646222530640399 1 0.0003651220530640399 1 0.0003651222530640399 1 0.0003656220530640399 1 0.0003656222530640399 1 0.0003661220530640399 1 0.0003661222530640399 1 0.0003666220530640399 1 0.0003666222530640399 1 0.0003671220530640399 1 0.00036712225306403994 1 0.00036732924646941807 1 0.0003673294464694181 1 0.0003725365334006625 1 0.0003725367334006625 1 0.0003728292464694181 1 0.0003728294464694181 1 0.0003733292464694181 1 0.0003733294464694181 1 0.0003738292464694181 1 0.00037382944646941813 1 0.00037432924646941813 1 0.00037432944646941814 1 0.00037482924646941814 1 0.00037482944646941816 1 0.00037532924646941816 1 0.00037532944646941817 1 0.00037582924646941817 1 0.0003758294464694182 1 0.0003763292464694182 1 0.0003763294464694182 1 0.0003768292464694182 1 0.0003768294464694182 1 0.0003773292464694182 1 0.0003773294464694182 1 0.0003775365334006625 1 0.0003775367334006625 1 0.00038274395561190434 1 0.00038274415561190435 1 0.0003830365334006625 1 0.00038303673340066253 1 0.0003835365334006625 1 0.0003835367334006625 1 0.00038403653340066243 1 0.00038403673340066245 1 0.0003845365334006624 1 0.0003845367334006624 1 0.00038503653340066235 1 0.00038503673340066236 1 0.0003855365334006623 1 0.0003855367334006623 1 0.00038603653340066226 1 0.0003860367334006623 1 0.0003865365334006622 1 0.00038653673340066224 1 0.0003870365334006622 1 0.0003870367334006622 1 0.00038753653340066214 1 0.00038753673340066215 1 0.0003877439556119038 1 0.0003877441556119038 1 0.00039295175422431375 1 0.00039295195422431377 1 0.00039324395561190383 1 0.00039324415561190385 1 0.00039374395561190384 1 0.00039374415561190386 1 0.00039424395561190386 1 0.00039424415561190387 1 0.00039474395561190387 1 0.0003947441556119039 1 0.0003952439556119039 1 0.0003952441556119039 1 0.0003957439556119039 1 0.0003957441556119039 1 0.0003962439556119039 1 0.0003962441556119039 1 0.0003967439556119039 1 0.00039674415561190393 1 0.00039724395561190393 1 0.00039724415561190394 1 0.00039774395561190394 1 0.00039774415561190396 1 0.00039795175422431377 1 0.0003979519542243138 1 0.00040315970887468036 1 0.00040315990887468037 1 0.00040345175422431385 1 0.00040345195422431386 1 0.0004039517542243139 1 0.0004039519542243139 1 0.000404451754224314 1 0.000404451954224314 1 0.00040495175422431405 1 0.00040495195422431406 1 0.0004054517542243141 1 0.0004054519542243141 1 0.0004059517542243142 1 0.0004059519542243142 1 0.00040645175422431424 1 0.00040645195422431426 1 0.0004069517542243143 1 0.0004069519542243143 1 0.0004074517542243144 1 0.0004074519542243144 1 0.00040795175422431444 1 0.00040795195422431446 1 0.0004081597088746809 1 0.0004081599088746809 1 0.0004133678210077549 1 0.0004133680210077549 1 0.0004136597088746809 1 0.0004136599088746809 1 0.00041415970887468095 1 0.00041415990887468096 1 0.000414659708874681 1 0.00041465990887468103 1 0.0004151597088746811 1 0.0004151599088746811 1 0.00041565970887468115 1 0.00041565990887468116 1 0.0004161597088746812 1 0.00041615990887468123 1 0.0004166597088746813 1 0.0004166599088746813 1 0.00041715970887468135 1 0.00041715990887468136 1 0.0004176597088746814 1 0.00041765990887468143 1 0.0004181597088746815 1 0.0004181599088746815 1 0.0004183678210077554 1 0.0004183680210077554 1 0.00042357605238244213 1 0.00042357625238244215 1 0.0004238678210077554 1 0.0004238680210077554 1 0.0004243678210077554 1 0.00042436802100775543 1 0.00042486782100775543 1 0.00042486802100775544 1 0.00042536782100775544 1 0.00042536802100775546 1 0.00042586782100775545 1 0.00042586802100775547 1 0.00042636782100775547 1 0.0004263680210077555 1 0.0004268678210077555 1 0.0004268680210077555 1 0.0004273678210077555 1 0.0004273680210077555 1 0.0004278678210077555 1 0.0004278680210077555 1 0.0004283678210077555 1 0.00042836802100775553 1 0.00042857605238244215 1 0.00042857625238244216 1 0.0004337845821168645 1 0.00043378478211686454 1 0.00043407605238244217 1 0.0004340762523824422 1 0.00043457605238244224 1 0.00043457625238244225 1 0.0004350760523824423 1 0.0004350762523824423 1 0.00043557605238244237 1 0.0004355762523824424 1 0.00043607605238244244 1 0.00043607625238244245 1 0.0004365760523824425 1 0.0004365762523824425 1 0.00043707605238244257 1 0.0004370762523824426 1 0.00043757605238244263 1 0.00043757625238244265 1 0.0004380760523824427 1 0.0004380762523824427 1 0.00043857605238244277 1 0.0004385762523824428 1 0.000438784582116865 1 0.00043878478211686504 1 0.00044399329473837737 1 0.0004439934947383774 1 0.00044428458211686505 1 0.00044428478211686506 1 0.00044478458211686506 1 0.0004447847821168651 1 0.0004452845821168651 1 0.0004452847821168651 1 0.0004457845821168651 1 0.0004457847821168651 1 0.0004462845821168651 1 0.0004462847821168651 1 0.0004467845821168651 1 0.0004467847821168651 1 0.0004472845821168651 1 0.00044728478211686514 1 0.00044778458211686514 1 0.00044778478211686515 1 0.00044828458211686515 1 0.00044828478211686516 1 0.00044878458211686516 1 0.0004487847821168652 1 0.0004489932947383774 1 0.0004489934947383774 1 0.0004542021916109949 1 0.0004542023916109949 1 0.0004544932947383774 1 0.0004544934947383774 1 0.00045499329473837737 1 0.0004549934947383774 1 0.0004554932947383773 1 0.00045549349473837734 1 0.0004559932947383773 1 0.0004559934947383773 1 0.00045649329473837724 1 0.00045649349473837725 1 0.0004569932947383772 1 0.0004569934947383772 1 0.00045749329473837716 1 0.00045749349473837717 1 0.0004579932947383771 1 0.00045799349473837713 1 0.00045849329473837707 1 0.0004584934947383771 1 0.00045899329473837703 1 0.00045899349473837704 1 0.00045920219161099435 1 0.00045920239161099436 1 0.00046441127816508496 1 0.00046441147816508497 1 0.0004647021916109944 1 0.0004647023916109944 1 0.0004652021916109944 1 0.0004652023916109944 1 0.0004657021916109944 1 0.0004657023916109944 1 0.0004662021916109944 1 0.0004662023916109944 1 0.0004667021916109944 1 0.00046670239161099444 1 0.00046720219161099444 1 0.00046720239161099445 1 0.00046770219161099445 1 0.00046770239161099446 1 0.00046820219161099446 1 0.0004682023916109945 1 0.00046870219161099447 1 0.0004687023916109945 1 0.0004692021916109945 1 0.0004692023916109945 1 0.00046941127816508497 1 0.000469411478165085 1 0.0004746205704165872 1 0.0004746207704165872 1 0.000474911278165085 1 0.000474911478165085 1 0.00047541127816508506 1 0.0004754114781650851 1 0.0004759112781650851 1 0.00047591147816508514 1 0.0004764112781650852 1 0.0004764114781650852 1 0.00047691127816508526 1 0.0004769114781650853 1 0.0004774112781650853 1 0.00047741147816508534 1 0.0004779112781650854 1 0.0004779114781650854 1 0.00047841127816508546 1 0.00047841147816508547 1 0.0004789112781650855 1 0.00047891147816508554 1 0.00047941127816508554 1 0.00047941147816508555 1 0.00047962057041658765 1 0.00047962077041658767 1 0.00048483012515769053 1 0.00048483032515769055 1 0.0004851205704165877 1 0.0004851207704165877 1 0.0004856205704165877 1 0.0004856207704165877 1 0.0004861205704165877 1 0.0004861207704165877 1 0.0004866205704165877 1 0.00048662077041658773 1 0.00048712057041658773 1 0.00048712077041658774 1 0.00048762057041658774 1 0.00048762077041658775 1 0.00048812057041658775 1 0.00048812077041658777 1 0.0004886205704165877 1 0.0004886207704165877 1 0.0004891205704165878 1 0.0004891207704165877 1 0.0004896205704165878 1 0.0004896207704165878 1 0.0004898301251576905 1 0.0004898303251576905 1 0.000495039780822236 1 0.000495039980822236 1 0.0004953301251576906 1 0.0004953303251576906 1 0.0004958301251576906 1 0.0004958303251576905 1 0.0004963301251576906 1 0.0004963303251576906 1 0.0004968301251576907 1 0.0004968303251576907 1 0.0004973301251576908 1 0.0004973303251576907 1 0.0004978301251576908 1 0.0004978303251576908 1 0.0004983301251576909 1 0.0004983303251576909 1 0.000498830125157691 1 0.0004988303251576909 1 0.000499330125157691 1 0.000499330325157691 1 0.0004998301251576911 1 0.0004998303251576911 1 0.0005000397808222364 1 0.0005000399808222363 1 0.0005052496159810823 1 0.0005052498159810822 1 0.0005055397808222363 1 0.0005055399808222363 1 0.0005060397808222364 1 0.0005060399808222364 1 0.0005065397808222365 1 0.0005065399808222364 1 0.0005070397808222365 1 0.0005070399808222365 1 0.0005075397808222366 1 0.0005075399808222366 1 0.0005080397808222367 1 0.0005080399808222366 1 0.0005085397808222367 1 0.0005085399808222367 1 0.0005090397808222368 1 0.0005090399808222368 1 0.0005095397808222369 1 0.0005095399808222368 1 0.000510039780822237 1 0.0005100399808222369 1 0.0005102496159810827 1)
X5 __ph_in[1]_v ph_in[1] __ph_in[1]_s 0 inout_sw_mod
V6 __ph_in[1]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 0 5.700184028257943e-06 0 5.7003840282579425e-06 1 6.200184028257943e-06 1 6.200384028257943e-06 0 6.700184028257943e-06 0 6.700384028257942e-06 1 7.200184028257943e-06 1 7.2003840282579425e-06 0 7.700184028257943e-06 0 7.700384028257944e-06 1 8.200184028257943e-06 1 8.200384028257944e-06 0 8.700184028257944e-06 0 8.700384028257944e-06 1 9.200184028257944e-06 1 9.200384028257945e-06 0 9.700184028257946e-06 0 9.700384028257947e-06 1 1.0200184028257948e-05 1 1.0200384028257949e-05 0 1.0400399910590747e-05 0 1.0400599910590748e-05 0 1.5900399910590747e-05 0 1.5900599910590748e-05 1 1.6400399910590746e-05 1 1.6400599910590746e-05 0 1.6900399910590744e-05 0 1.6900599910590745e-05 1 1.7400399910590743e-05 1 1.7400599910590743e-05 0 1.790039991059074e-05 0 1.7900599910590742e-05 1 1.840039991059074e-05 1 1.840059991059074e-05 0 1.890039991059074e-05 0 1.890059991059074e-05 1 1.9400399910590737e-05 1 1.9400599910590738e-05 0 1.9900399910590736e-05 0 1.9900599910590736e-05 1 2.0400399910590735e-05 1 2.0400599910590735e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 0 2.6100911580126336e-05 0 2.6101111580126337e-05 1 2.6600911580126335e-05 1 2.6601111580126335e-05 0 2.7100911580126333e-05 0 2.7101111580126334e-05 1 2.7600911580126332e-05 1 2.7601111580126332e-05 0 2.810091158012633e-05 0 2.810111158012633e-05 1 2.860091158012633e-05 1 2.860111158012633e-05 0 2.9100911580126328e-05 0 2.9101111580126328e-05 1 2.9600911580126326e-05 1 2.9601111580126327e-05 0 3.0100911580126325e-05 0 3.0101111580126325e-05 1 3.0600911580126324e-05 1 3.0601111580126324e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 0 3.630158374751402e-05 0 3.630178374751402e-05 1 3.680158374751402e-05 1 3.680178374751402e-05 0 3.730158374751402e-05 0 3.730178374751402e-05 1 3.780158374751402e-05 1 3.780178374751402e-05 0 3.8301583747514016e-05 0 3.8301783747514016e-05 1 3.8801583747514014e-05 1 3.8801783747514015e-05 0 3.930158374751401e-05 0 3.9301783747514013e-05 1 3.980158374751401e-05 1 3.980178374751401e-05 0 4.030158374751401e-05 0 4.030178374751401e-05 1 4.080158374751401e-05 1 4.080178374751401e-05 0 4.1002390731437404e-05 0 4.1002590731437404e-05 0 4.65023907314374e-05 0 4.65025907314374e-05 1 4.70023907314374e-05 1 4.70025907314374e-05 0 4.75023907314374e-05 0 4.75025907314374e-05 1 4.80023907314374e-05 1 4.80025907314374e-05 0 4.8502390731437396e-05 0 4.85025907314374e-05 1 4.9002390731437395e-05 1 4.9002590731437395e-05 0 4.9502390731437394e-05 0 4.9502590731437394e-05 1 5.000239073143739e-05 1 5.000259073143739e-05 0 5.050239073143739e-05 0 5.050259073143739e-05 1 5.100239073143739e-05 1 5.100259073143739e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 0 5.670345687967774e-05 0 5.670365687967774e-05 1 5.720345687967774e-05 1 5.720365687967774e-05 0 5.770345687967774e-05 0 5.770365687967774e-05 1 5.820345687967774e-05 1 5.820365687967774e-05 0 5.870345687967774e-05 0 5.870365687967774e-05 1 5.9203456879677736e-05 1 5.9203656879677736e-05 0 5.9703456879677734e-05 0 5.9703656879677735e-05 1 6.020345687967773e-05 1 6.020365687967773e-05 0 6.070345687967773e-05 0 6.070365687967773e-05 1 6.120345687967773e-05 1 6.120365687967773e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 0 6.690480297716098e-05 0 6.690500297716098e-05 1 6.740480297716097e-05 1 6.740500297716097e-05 0 6.790480297716095e-05 0 6.790500297716095e-05 1 6.840480297716094e-05 1 6.840500297716094e-05 0 6.890480297716092e-05 0 6.890500297716092e-05 1 6.94048029771609e-05 1 6.940500297716091e-05 0 6.990480297716089e-05 0 6.990500297716089e-05 1 7.040480297716088e-05 1 7.040500297716088e-05 0 7.090480297716086e-05 0 7.090500297716086e-05 1 7.140480297716085e-05 1 7.140500297716085e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 0 7.710630340083568e-05 0 7.710650340083568e-05 1 7.760630340083568e-05 1 7.760650340083568e-05 0 7.810630340083568e-05 0 7.810650340083568e-05 1 7.860630340083568e-05 1 7.860650340083568e-05 0 7.910630340083568e-05 0 7.910650340083568e-05 1 7.960630340083567e-05 1 7.960650340083567e-05 0 8.010630340083567e-05 0 8.010650340083567e-05 1 8.060630340083567e-05 1 8.060650340083567e-05 0 8.110630340083567e-05 0 8.110650340083567e-05 1 8.160630340083567e-05 1 8.160650340083567e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 0 8.73080003149639e-05 0 8.73082003149639e-05 1 8.780800031496389e-05 1 8.780820031496389e-05 0 8.830800031496387e-05 0 8.830820031496387e-05 1 8.880800031496386e-05 1 8.880820031496386e-05 0 8.930800031496384e-05 0 8.930820031496384e-05 1 8.980800031496383e-05 1 8.980820031496383e-05 0 9.030800031496381e-05 0 9.030820031496381e-05 1 9.08080003149638e-05 1 9.08082003149638e-05 0 9.130800031496378e-05 0 9.130820031496378e-05 1 9.180800031496377e-05 1 9.180820031496377e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 0 9.750984556640299e-05 0 9.751004556640299e-05 1 9.8009845566403e-05 1 9.8010045566403e-05 0 9.850984556640302e-05 0 9.851004556640302e-05 1 9.900984556640303e-05 1 9.901004556640303e-05 0 9.950984556640304e-05 0 9.951004556640304e-05 1 0.00010000984556640305 1 0.00010001004556640305 0 0.00010050984556640307 0 0.00010051004556640307 1 0.00010100984556640308 1 0.00010101004556640308 0 0.00010150984556640309 0 0.00010151004556640309 1 0.0001020098455664031 1 0.0001020100455664031 0 0.00010221189158154771 0 0.00010221209158154771 0 0.00010771189158154771 0 0.00010771209158154771 1 0.0001082118915815477 1 0.0001082120915815477 0 0.00010871189158154768 0 0.00010871209158154768 1 0.00010921189158154767 1 0.00010921209158154767 0 0.00010971189158154765 0 0.00010971209158154765 1 0.00011021189158154764 1 0.00011021209158154764 0 0.00011071189158154762 0 0.00011071209158154762 1 0.00011121189158154761 1 0.00011121209158154761 0 0.00011171189158154759 0 0.00011171209158154759 1 0.00011221189158154758 1 0.00011221209158154758 0 0.00011241412374722472 0 0.00011241432374722472 0 0.0001179141237472247 0 0.0001179143237472247 1 0.00011841412374722469 1 0.00011841432374722469 0 0.00011891412374722467 0 0.00011891432374722467 1 0.00011941412374722466 1 0.00011941432374722466 0 0.00011991412374722464 0 0.00011991432374722464 1 0.00012041412374722463 1 0.00012041432374722463 0 0.00012091412374722461 0 0.00012091432374722461 1 0.00012141412374722461 1 0.00012141432374722461 0 0.00012191412374722461 0 0.00012191432374722461 1 0.0001224141237472246 1 0.00012241432374722458 0 0.00012261667966227715 0 0.00012261687966227714 0 0.00012811667966227717 0 0.00012811687966227716 1 0.00012861667966227719 1 0.00012861687966227717 0 0.0001291166796622772 0 0.00012911687966227719 1 0.0001296166796622772 1 0.0001296168796622772 0 0.00013011667966227722 0 0.0001301168796622772 1 0.00013061667966227723 1 0.00013061687966227722 0 0.00013111667966227725 0 0.00013111687966227723 1 0.00013161667966227726 1 0.00013161687966227725 0 0.00013211667966227727 0 0.00013211687966227726 1 0.00013261667966227728 1 0.00013261687966227727 0 0.00013281929267817236 0 0.00013281949267817235 0 0.0001383192926781724 0 0.00013831949267817238 1 0.0001388192926781724 1 0.0001388194926781724 0 0.00013931929267817241 0 0.0001393194926781724 1 0.00013981929267817243 1 0.0001398194926781724 0 0.00014031929267817244 0 0.00014031949267817242 1 0.00014081929267817245 1 0.00014081949267817244 0 0.00014131929267817246 0 0.00014131949267817245 1 0.00014181929267817247 1 0.00014181949267817246 0 0.0001423192926781725 0 0.00014231949267817247 1 0.0001428192926781725 1 0.00014281949267817249 0 0.00014302214851901298 0 0.00014302234851901297 0 0.000148522148519013 0 0.000148522348519013 1 0.00014902214851901302 1 0.000149022348519013 0 0.00014952214851901303 0 0.00014952234851901302 1 0.00015002214851901304 1 0.00015002234851901303 0 0.00015052214851901305 0 0.00015052234851901304 1 0.00015102214851901307 1 0.00015102234851901305 0 0.00015152214851901308 0 0.00015152234851901306 1 0.0001520221485190131 1 0.00015202234851901308 0 0.0001525221485190131 0 0.0001525223485190131 1 0.00015302214851901311 1 0.0001530223485190131 0 0.00015322531083256498 0 0.00015322551083256497 0 0.000158725310832565 0 0.000158725510832565 1 0.00015922531083256502 1 0.000159225510832565 0 0.00015972531083256503 0 0.00015972551083256502 1 0.00016022531083256504 1 0.00016022551083256503 0 0.00016072531083256505 0 0.00016072551083256504 1 0.00016122531083256507 1 0.00016122551083256505 0 0.00016172531083256508 0 0.00016172551083256506 1 0.0001622253108325651 1 0.00016222551083256508 0 0.0001627253108325651 0 0.0001627255108325651 1 0.00016322531083256511 1 0.0001632255108325651 0 0.0001634286310398012 0 0.00016342883103980118 0 0.0001689286310398012 0 0.00016892883103980118 1 0.0001694286310398012 1 0.0001694288310398012 0 0.00016992863103980121 0 0.0001699288310398012 1 0.00017042863103980123 1 0.0001704288310398012 0 0.00017092863103980124 0 0.00017092883103980122 1 0.00017142863103980125 1 0.00017142883103980124 0 0.00017192863103980126 0 0.00017192883103980125 1 0.00017242863103980127 1 0.00017242883103980126 0 0.0001729286310398013 0 0.00017292883103980127 1 0.0001734286310398013 1 0.00017342883103980129 0 0.0001736321391540218 0 0.0001736323391540218 0 0.00017913213915402183 0 0.00017913233915402182 1 0.00017963213915402185 1 0.00017963233915402183 0 0.00018013213915402186 0 0.00018013233915402185 1 0.00018063213915402187 1 0.00018063233915402186 0 0.00018113213915402188 0 0.00018113233915402187 1 0.0001816321391540219 1 0.00018163233915402188 0 0.0001821321391540219 0 0.0001821323391540219 1 0.00018263213915402192 1 0.0001826323391540219 0 0.00018313213915402193 0 0.00018313233915402192 1 0.00018363213915402194 1 0.00018363233915402193 0 0.0001838358186013159 0 0.00018383601860131587 0 0.0001893358186013159 0 0.0001893360186013159 1 0.00018983581860131592 1 0.0001898360186013159 0 0.00019033581860131594 0 0.00019033601860131592 1 0.00019083581860131595 1 0.00019083601860131594 0 0.00019133581860131596 0 0.00019133601860131595 1 0.00019183581860131597 1 0.00019183601860131596 0 0.00019233581860131599 0 0.00019233601860131597 1 0.000192835818601316 1 0.00019283601860131598 0 0.000193335818601316 0 0.000193336018601316 1 0.00019383581860131602 1 0.000193836018601316 0 0.00019403971249211136 0 0.00019403991249211135 0 0.00019953971249211139 0 0.00019953991249211137 1 0.0002000397124921114 1 0.00020003991249211139 0 0.0002005397124921114 0 0.0002005399124921114 1 0.00020103971249211142 1 0.0002010399124921114 0 0.00020153971249211143 0 0.00020153991249211142 1 0.00020203971249211145 1 0.00020203991249211143 0 0.00020253971249211146 0 0.00020253991249211145 1 0.00020303971249211147 1 0.00020303991249211146 0 0.00020353971249211148 0 0.00020353991249211147 1 0.0002040397124921115 1 0.00020403991249211148 0 0.0002042437273079041 0 0.00020424392730790408 0 0.00020974372730790412 0 0.0002097439273079041 1 0.00021024372730790413 1 0.00021024392730790412 0 0.00021074372730790414 0 0.00021074392730790413 1 0.00021124372730790415 1 0.00021124392730790414 0 0.00021174372730790416 0 0.00021174392730790415 1 0.00021224372730790418 1 0.00021224392730790416 0 0.0002127437273079042 0 0.00021274392730790418 1 0.0002132437273079042 1 0.0002132439273079042 0 0.0002137437273079042 0 0.0002137439273079042 1 0.00021424372730790423 1 0.0002142439273079042 0 0.00021444808721675775 0 0.00021444828721675773 0 0.00021994808721675777 0 0.00021994828721675776 1 0.00022044808721675778 1 0.00022044828721675777 0 0.0002209480872167578 0 0.00022094828721675778 1 0.0002214480872167578 1 0.0002214482872167578 0 0.00022194808721675782 0 0.0002219482872167578 1 0.00022244808721675783 1 0.00022244828721675782 0 0.00022294808721675784 0 0.00022294828721675783 1 0.00022344808721675786 1 0.00022344828721675784 0 0.00022394808721675787 0 0.00022394828721675786 1 0.00022444808721675788 1 0.00022444828721675787 0 0.00022465261116331255 0 0.00022465281116331253 0 0.00023015261116331257 0 0.00023015281116331256 1 0.00023065261116331259 1 0.00023065281116331257 0 0.0002311526111633126 0 0.00023115281116331258 1 0.0002316526111633126 1 0.0002316528111633126 0 0.00023215261116331262 0 0.0002321528111633126 1 0.00023265261116331263 1 0.00023265281116331262 0 0.00023315261116331265 0 0.00023315281116331263 1 0.00023365261116331266 1 0.00023365281116331265 0 0.00023415261116331267 0 0.00023415281116331266 1 0.00023465261116331268 1 0.00023465281116331267 0 0.00023485725348777872 0 0.0002348574534877787 0 0.00024035725348777874 0 0.00024035745348777873 1 0.00024085725348777876 1 0.00024085745348777874 0 0.00024135725348777877 0 0.00024135745348777876 1 0.00024185725348777878 1 0.00024185745348777877 0 0.0002423572534877788 0 0.00024235745348777878 1 0.0002428572534877788 1 0.0002428574534877788 0 0.00024335725348777882 0 0.0002433574534877788 1 0.00024385725348777883 1 0.00024385745348777882 0 0.00024435725348777884 0 0.00024435745348777886 1 0.0002448572534877788 1 0.0002448574534877788 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025056213249421646 0 0.0002505623324942165 1 0.0002510621324942165 1 0.0002510623324942165 0 0.0002515621324942165 0 0.0002515623324942165 1 0.0002520621324942165 1 0.0002520623324942165 0 0.0002525621324942165 0 0.0002525623324942165 1 0.0002530621324942165 1 0.00025306233249421654 0 0.00025356213249421654 0 0.00025356233249421655 1 0.00025406213249421655 1 0.00025406233249421656 0 0.00025456213249421656 0 0.0002545623324942166 1 0.00025506213249421646 1 0.0002550623324942165 0 0.00025526732409400483 0 0.00025526752409400484 0 0.00026076732409400485 0 0.00026076752409400487 1 0.0002612673240940049 1 0.00026126752409400493 0 0.000261767324094005 0 0.000261767524094005 1 0.00026226732409400505 1 0.00026226752409400507 0 0.0002627673240940051 0 0.00026276752409400513 1 0.0002632673240940052 1 0.0002632675240940052 0 0.00026376732409400525 0 0.00026376752409400527 1 0.0002642673240940053 1 0.00026426752409400533 0 0.0002647673240940054 0 0.0002647675240940054 1 0.00026526732409400534 1 0.00026526752409400536 0 0.0002654725372742233 0 0.00026547273727422333 0 0.00027097253727422334 0 0.00027097273727422336 1 0.0002714725372742233 1 0.0002714727372742233 0 0.00027197253727422326 0 0.00027197273727422327 1 0.0002724725372742232 1 0.00027247273727422323 0 0.0002729725372742232 0 0.0002729727372742232 1 0.00027347253727422313 1 0.00027347273727422315 0 0.0002739725372742231 0 0.0002739727372742231 1 0.00027447253727422305 1 0.00027447273727422306 0 0.000274972537274223 0 0.000274972737274223 1 0.00027547253727422285 1 0.00027547273727422287 0 0.0002756781009094726 0 0.0002756783009094726 0 0.0002811781009094726 0 0.0002811783009094726 1 0.0002816781009094726 1 0.00028167830090947263 0 0.0002821781009094726 0 0.00028217830090947264 1 0.00028267810090947264 1 0.00028267830090947265 0 0.00028317810090947265 0 0.00028317830090947266 1 0.00028367810090947266 1 0.0002836783009094727 0 0.0002841781009094727 0 0.0002841783009094727 1 0.0002846781009094727 1 0.0002846783009094727 0 0.0002851781009094727 0 0.0002851783009094727 1 0.0002856781009094726 1 0.0002856783009094726 0 0.0002858838383549405 0 0.0002858840383549405 0 0.00029138383835494047 0 0.0002913840383549405 1 0.0002918838383549404 1 0.00029188403835494044 0 0.0002923838383549404 0 0.0002923840383549404 1 0.00029288383835494034 1 0.00029288403835494035 0 0.0002933838383549403 0 0.0002933840383549403 1 0.00029388383835494026 1 0.00029388403835494027 0 0.0002943838383549402 0 0.00029438403835494023 1 0.00029488383835494017 1 0.0002948840383549402 0 0.00029538383835494013 0 0.00029538403835494014 1 0.00029588383835494 1 0.00029588403835494 0 0.0002960896923277906 0 0.00029608989232779063 0 0.0003015896923277906 0 0.0003015898923277906 1 0.00030208969232779054 1 0.00030208989232779056 0 0.0003025896923277905 0 0.0003025898923277905 1 0.00030308969232779046 1 0.00030308989232779047 0 0.0003035896923277904 0 0.00030358989232779043 1 0.0003040896923277904 1 0.0003040898923277904 0 0.00030458969232779033 0 0.00030458989232779035 1 0.0003050896923277903 1 0.0003050898923277903 0 0.00030558969232779025 0 0.00030558989232779026 1 0.0003060896923277901 1 0.0003060898923277901 0 0.0003062957259554461 0 0.0003062959259554461 0 0.00031179572595544606 0 0.00031179592595544607 1 0.000312295725955446 1 0.00031229592595544603 0 0.000312795725955446 0 0.000312795925955446 1 0.00031329572595544593 1 0.00031329592595544595 0 0.0003137957259554459 0 0.0003137959259554459 1 0.00031429572595544585 1 0.00031429592595544586 0 0.0003147957259554458 0 0.0003147959259554458 1 0.00031529572595544576 1 0.0003152959259554458 0 0.0003157957259554457 0 0.00031579592595544574 1 0.00031629572595544557 1 0.0003162959259554456 0 0.0003165020377403174 0 0.0003165022377403174 0 0.00032200203774031743 0 0.00032200223774031745 1 0.0003225020377403175 1 0.0003225022377403175 0 0.00032300203774031757 0 0.0003230022377403176 1 0.00032350203774031763 1 0.00032350223774031765 0 0.0003240020377403177 0 0.0003240022377403177 1 0.00032450203774031777 1 0.0003245022377403178 0 0.00032500203774031783 0 0.00032500223774031785 1 0.0003255020377403179 1 0.0003255022377403179 0 0.00032600203774031796 0 0.000326002237740318 1 0.0003265020377403179 1 0.00032650223774031794 0 0.0003267084673472993 0 0.0003267086673472993 0 0.0003322084673472994 0 0.0003322086673472994 1 0.00033270846734729945 1 0.00033270866734729946 0 0.0003332084673472995 0 0.00033320866734729953 1 0.0003337084673472996 1 0.0003337086673472996 0 0.00033420846734729965 0 0.00033420866734729966 1 0.0003347084673472997 1 0.00033470866734729973 0 0.0003352084673472998 0 0.0003352086673472998 1 0.00033570846734729985 1 0.00033570866734729986 0 0.0003362084673472999 0 0.00033620866734729993 1 0.00033670846734729987 1 0.0003367086673472999 0 0.00033691523365255696 0 0.000336915433652557 0 0.00034241523365255693 0 0.00034241543365255695 1 0.0003429152336525569 1 0.0003429154336525569 0 0.00034341523365255685 0 0.00034341543365255686 1 0.0003439152336525568 1 0.0003439154336525568 0 0.00034441523365255676 0 0.0003444154336525568 1 0.0003449152336525567 1 0.00034491543365255674 0 0.0003454152336525567 0 0.0003454154336525567 1 0.00034591523365255664 1 0.00034591543365255665 0 0.0003464152336525566 0 0.0003464154336525566 1 0.00034691523365255644 1 0.00034691543365255646 0 0.00034712205306404025 0 0.00034712225306404026 0 0.0003526220530640403 0 0.0003526222530640403 1 0.00035312205306404023 1 0.00035312225306404025 0 0.0003536220530640402 0 0.0003536222530640402 1 0.00035412205306404015 1 0.00035412225306404016 0 0.0003546220530640401 0 0.0003546222530640401 1 0.00035512205306404007 1 0.0003551222530640401 0 0.00035562205306404 0 0.00035562225306404004 1 0.00035612205306404 1 0.00035612225306404 0 0.00035662205306403994 0 0.00035662225306403995 1 0.0003571220530640398 1 0.0003571222530640398 0 0.00035732924646941804 0 0.00035732944646941806 0 0.00036282924646941807 0 0.0003628294464694181 1 0.0003633292464694181 1 0.0003633294464694181 0 0.0003638292464694181 0 0.0003638294464694181 1 0.0003643292464694181 1 0.0003643294464694181 0 0.0003648292464694181 0 0.00036482944646941813 1 0.00036532924646941813 1 0.00036532944646941814 0 0.00036582924646941814 0 0.00036582944646941815 1 0.00036632924646941815 1 0.00036632944646941817 0 0.00036682924646941817 0 0.0003668294464694182 1 0.00036732924646941807 1 0.0003673294464694181 0 0.00036753653340066246 0 0.0003675367334006625 0 0.0003730365334006625 0 0.0003730367334006625 1 0.0003735365334006625 1 0.0003735367334006625 0 0.0003740365334006625 0 0.00037403673340066253 1 0.0003745365334006625 1 0.00037453673340066254 0 0.00037503653340066254 0 0.00037503673340066255 1 0.00037553653340066255 1 0.00037553673340066256 0 0.00037603653340066256 0 0.0003760367334006626 1 0.0003765365334006626 1 0.0003765367334006626 0 0.0003770365334006626 0 0.0003770367334006626 1 0.0003775365334006625 1 0.0003775367334006625 0 0.0003777439556119043 0 0.00037774415561190434 0 0.0003832439556119043 0 0.0003832441556119043 1 0.00038374395561190425 1 0.00038374415561190427 0 0.0003842439556119042 0 0.0003842441556119042 1 0.00038474395561190417 1 0.0003847441556119042 0 0.0003852439556119041 0 0.00038524415561190414 1 0.0003857439556119041 1 0.0003857441556119041 0 0.00038624395561190404 0 0.00038624415561190406 1 0.000386743955611904 1 0.000386744155611904 0 0.00038724395561190396 0 0.00038724415561190397 1 0.0003877439556119038 1 0.0003877441556119038 0 0.00038795175422431374 0 0.00038795195422431375 0 0.00039345175422431377 0 0.0003934519542243138 1 0.0003939517542243138 1 0.0003939519542243138 0 0.0003944517542243138 0 0.0003944519542243138 1 0.0003949517542243138 1 0.0003949519542243138 0 0.0003954517542243138 0 0.00039545195422431383 1 0.0003959517542243138 1 0.00039595195422431384 0 0.00039645175422431384 0 0.00039645195422431385 1 0.00039695175422431385 1 0.00039695195422431386 0 0.00039745175422431386 0 0.0003974519542243139 1 0.00039795175422431377 1 0.0003979519542243138 0 0.00039815970887468034 0 0.00039815990887468036 0 0.0004036597088746804 0 0.00040365990887468044 1 0.0004041597088746805 1 0.0004041599088746805 0 0.00040465970887468056 0 0.00040465990887468057 1 0.0004051597088746806 1 0.00040515990887468064 0 0.0004056597088746807 0 0.0004056599088746807 1 0.00040615970887468076 1 0.00040615990887468077 0 0.0004066597088746808 0 0.00040665990887468084 1 0.0004071597088746809 1 0.0004071599088746809 0 0.00040765970887468095 0 0.00040765990887468097 1 0.0004081597088746809 1 0.0004081599088746809 0 0.00040836782100775487 0 0.0004083680210077549 0 0.0004138678210077549 0 0.0004138680210077549 1 0.00041436782100775496 1 0.00041436802100775497 0 0.000414867821007755 0 0.00041486802100775504 1 0.0004153678210077551 1 0.0004153680210077551 0 0.00041586782100775516 0 0.00041586802100775517 1 0.0004163678210077552 1 0.00041636802100775524 0 0.0004168678210077553 0 0.0004168680210077553 1 0.00041736782100775536 1 0.00041736802100775537 0 0.0004178678210077554 0 0.00041786802100775544 1 0.0004183678210077554 1 0.0004183680210077554 0 0.0004185760523824421 0 0.00041857625238244213 0 0.00042407605238244214 0 0.00042407625238244216 1 0.00042457605238244216 1 0.00042457625238244217 0 0.00042507605238244217 0 0.0004250762523824422 1 0.0004255760523824422 1 0.0004255762523824422 0 0.0004260760523824422 0 0.0004260762523824422 1 0.0004265760523824422 1 0.0004265762523824422 0 0.0004270760523824422 0 0.00042707625238244223 1 0.00042757605238244223 1 0.00042757625238244224 0 0.00042807605238244224 0 0.00042807625238244226 1 0.00042857605238244215 1 0.00042857625238244216 0 0.0004287845821168645 0 0.0004287847821168645 0 0.00043428458211686454 0 0.00043428478211686455 1 0.0004347845821168646 1 0.0004347847821168646 0 0.00043528458211686467 0 0.0004352847821168647 1 0.00043578458211686474 1 0.00043578478211686475 0 0.0004362845821168648 0 0.0004362847821168648 1 0.00043678458211686487 1 0.0004367847821168649 0 0.00043728458211686493 0 0.00043728478211686495 1 0.000437784582116865 1 0.000437784782116865 0 0.00043828458211686507 0 0.0004382847821168651 1 0.000438784582116865 1 0.00043878478211686504 0 0.00043899329473837736 0 0.00043899349473837737 0 0.0004444932947383774 0 0.0004444934947383774 1 0.0004449932947383774 1 0.0004449934947383774 0 0.0004454932947383774 0 0.0004454934947383774 1 0.0004459932947383774 1 0.00044599349473837743 0 0.00044649329473837743 0 0.00044649349473837745 1 0.00044699329473837744 1 0.00044699349473837746 0 0.00044749329473837746 0 0.00044749349473837747 1 0.00044799329473837747 1 0.0004479934947383775 0 0.0004484932947383775 0 0.0004484934947383775 1 0.0004489932947383774 1 0.0004489934947383774 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045470219161099484 0 0.00045470239161099485 1 0.0004552021916109948 1 0.0004552023916109948 0 0.00045570219161099475 0 0.00045570239161099477 1 0.0004562021916109947 1 0.0004562023916109947 0 0.00045670219161099467 0 0.0004567023916109947 1 0.0004572021916109946 1 0.00045720239161099464 0 0.0004577021916109946 0 0.0004577023916109946 1 0.00045820219161099454 1 0.00045820239161099456 0 0.0004587021916109945 0 0.0004587023916109945 1 0.00045920219161099435 1 0.00045920239161099436 0 0.00045941127816508494 0 0.00045941147816508496 0 0.00046491127816508497 0 0.000464911478165085 1 0.000465411278165085 1 0.000465411478165085 0 0.000465911278165085 0 0.000465911478165085 1 0.000466411278165085 1 0.000466411478165085 0 0.000466911278165085 0 0.00046691147816508503 1 0.00046741127816508503 1 0.00046741147816508504 0 0.00046791127816508504 0 0.00046791147816508506 1 0.00046841127816508505 1 0.00046841147816508507 0 0.00046891127816508507 0 0.0004689114781650851 1 0.00046941127816508497 1 0.000469411478165085 0 0.0004696205704165872 0 0.0004696207704165872 0 0.0004751205704165872 0 0.00047512077041658723 1 0.0004756205704165873 1 0.0004756207704165873 0 0.00047612057041658735 0 0.00047612077041658737 1 0.0004766205704165874 1 0.00047662077041658743 0 0.0004771205704165875 0 0.0004771207704165875 1 0.00047762057041658755 1 0.00047762077041658757 0 0.0004781205704165876 0 0.00047812077041658763 1 0.0004786205704165877 1 0.0004786207704165877 0 0.00047912057041658775 0 0.00047912077041658776 1 0.00047962057041658765 1 0.00047962077041658767 0 0.0004798301251576905 0 0.00047983032515769053 0 0.00048533012515769054 0 0.00048533032515769056 1 0.00048583012515769056 1 0.00048583032515769057 0 0.00048633012515769057 0 0.0004863303251576906 1 0.0004868301251576906 1 0.0004868303251576906 0 0.0004873301251576906 0 0.0004873303251576906 1 0.0004878301251576906 1 0.0004878303251576906 0 0.0004883301251576906 0 0.0004883303251576905 1 0.0004888301251576906 1 0.0004888303251576906 0 0.0004893301251576907 0 0.0004893303251576907 1 0.0004898301251576905 1 0.0004898303251576905 0 0.000490039780822236 0 0.000490039980822236 0 0.000495539780822236 0 0.000495539980822236 1 0.0004960397808222361 1 0.000496039980822236 0 0.0004965397808222361 0 0.0004965399808222361 1 0.0004970397808222362 1 0.0004970399808222362 0 0.0004975397808222363 0 0.0004975399808222362 1 0.0004980397808222363 1 0.0004980399808222363 0 0.0004985397808222364 0 0.0004985399808222364 1 0.0004990397808222365 1 0.0004990399808222364 0 0.0004995397808222365 0 0.0004995399808222365 1 0.0005000397808222364 1 0.0005000399808222363 0 0.0005002496159810823 0 0.0005002498159810822 0 0.0005057496159810823 0 0.0005057498159810823 1 0.0005062496159810824 1 0.0005062498159810824 0 0.0005067496159810825 0 0.0005067498159810824 1 0.0005072496159810825 1 0.0005072498159810825 0 0.0005077496159810826 0 0.0005077498159810826 1 0.0005082496159810827 1 0.0005082498159810826 0 0.0005087496159810827 0 0.0005087498159810827 1 0.0005092496159810828 1 0.0005092498159810828 0 0.0005097496159810829 0 0.0005097498159810828 1 0.0005102496159810827 0)
V7 __ph_in[1]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 5.700184028257943e-06 1 5.7003840282579425e-06 1 6.200184028257943e-06 1 6.200384028257943e-06 1 6.700184028257943e-06 1 6.700384028257942e-06 1 7.200184028257943e-06 1 7.2003840282579425e-06 1 7.700184028257943e-06 1 7.700384028257944e-06 1 8.200184028257943e-06 1 8.200384028257944e-06 1 8.700184028257944e-06 1 8.700384028257944e-06 1 9.200184028257944e-06 1 9.200384028257945e-06 1 9.700184028257946e-06 1 9.700384028257947e-06 1 1.0200184028257948e-05 1 1.0200384028257949e-05 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 1.5900399910590747e-05 1 1.5900599910590748e-05 1 1.6400399910590746e-05 1 1.6400599910590746e-05 1 1.6900399910590744e-05 1 1.6900599910590745e-05 1 1.7400399910590743e-05 1 1.7400599910590743e-05 1 1.790039991059074e-05 1 1.7900599910590742e-05 1 1.840039991059074e-05 1 1.840059991059074e-05 1 1.890039991059074e-05 1 1.890059991059074e-05 1 1.9400399910590737e-05 1 1.9400599910590738e-05 1 1.9900399910590736e-05 1 1.9900599910590736e-05 1 2.0400399910590735e-05 1 2.0400599910590735e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 2.6100911580126336e-05 1 2.6101111580126337e-05 1 2.6600911580126335e-05 1 2.6601111580126335e-05 1 2.7100911580126333e-05 1 2.7101111580126334e-05 1 2.7600911580126332e-05 1 2.7601111580126332e-05 1 2.810091158012633e-05 1 2.810111158012633e-05 1 2.860091158012633e-05 1 2.860111158012633e-05 1 2.9100911580126328e-05 1 2.9101111580126328e-05 1 2.9600911580126326e-05 1 2.9601111580126327e-05 1 3.0100911580126325e-05 1 3.0101111580126325e-05 1 3.0600911580126324e-05 1 3.0601111580126324e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 3.630158374751402e-05 1 3.630178374751402e-05 1 3.680158374751402e-05 1 3.680178374751402e-05 1 3.730158374751402e-05 1 3.730178374751402e-05 1 3.780158374751402e-05 1 3.780178374751402e-05 1 3.8301583747514016e-05 1 3.8301783747514016e-05 1 3.8801583747514014e-05 1 3.8801783747514015e-05 1 3.930158374751401e-05 1 3.9301783747514013e-05 1 3.980158374751401e-05 1 3.980178374751401e-05 1 4.030158374751401e-05 1 4.030178374751401e-05 1 4.080158374751401e-05 1 4.080178374751401e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 4.65023907314374e-05 1 4.65025907314374e-05 1 4.70023907314374e-05 1 4.70025907314374e-05 1 4.75023907314374e-05 1 4.75025907314374e-05 1 4.80023907314374e-05 1 4.80025907314374e-05 1 4.8502390731437396e-05 1 4.85025907314374e-05 1 4.9002390731437395e-05 1 4.9002590731437395e-05 1 4.9502390731437394e-05 1 4.9502590731437394e-05 1 5.000239073143739e-05 1 5.000259073143739e-05 1 5.050239073143739e-05 1 5.050259073143739e-05 1 5.100239073143739e-05 1 5.100259073143739e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 5.670345687967774e-05 1 5.670365687967774e-05 1 5.720345687967774e-05 1 5.720365687967774e-05 1 5.770345687967774e-05 1 5.770365687967774e-05 1 5.820345687967774e-05 1 5.820365687967774e-05 1 5.870345687967774e-05 1 5.870365687967774e-05 1 5.9203456879677736e-05 1 5.9203656879677736e-05 1 5.9703456879677734e-05 1 5.9703656879677735e-05 1 6.020345687967773e-05 1 6.020365687967773e-05 1 6.070345687967773e-05 1 6.070365687967773e-05 1 6.120345687967773e-05 1 6.120365687967773e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 6.690480297716098e-05 1 6.690500297716098e-05 1 6.740480297716097e-05 1 6.740500297716097e-05 1 6.790480297716095e-05 1 6.790500297716095e-05 1 6.840480297716094e-05 1 6.840500297716094e-05 1 6.890480297716092e-05 1 6.890500297716092e-05 1 6.94048029771609e-05 1 6.940500297716091e-05 1 6.990480297716089e-05 1 6.990500297716089e-05 1 7.040480297716088e-05 1 7.040500297716088e-05 1 7.090480297716086e-05 1 7.090500297716086e-05 1 7.140480297716085e-05 1 7.140500297716085e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 7.710630340083568e-05 1 7.710650340083568e-05 1 7.760630340083568e-05 1 7.760650340083568e-05 1 7.810630340083568e-05 1 7.810650340083568e-05 1 7.860630340083568e-05 1 7.860650340083568e-05 1 7.910630340083568e-05 1 7.910650340083568e-05 1 7.960630340083567e-05 1 7.960650340083567e-05 1 8.010630340083567e-05 1 8.010650340083567e-05 1 8.060630340083567e-05 1 8.060650340083567e-05 1 8.110630340083567e-05 1 8.110650340083567e-05 1 8.160630340083567e-05 1 8.160650340083567e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 8.73080003149639e-05 1 8.73082003149639e-05 1 8.780800031496389e-05 1 8.780820031496389e-05 1 8.830800031496387e-05 1 8.830820031496387e-05 1 8.880800031496386e-05 1 8.880820031496386e-05 1 8.930800031496384e-05 1 8.930820031496384e-05 1 8.980800031496383e-05 1 8.980820031496383e-05 1 9.030800031496381e-05 1 9.030820031496381e-05 1 9.08080003149638e-05 1 9.08082003149638e-05 1 9.130800031496378e-05 1 9.130820031496378e-05 1 9.180800031496377e-05 1 9.180820031496377e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 9.750984556640299e-05 1 9.751004556640299e-05 1 9.8009845566403e-05 1 9.8010045566403e-05 1 9.850984556640302e-05 1 9.851004556640302e-05 1 9.900984556640303e-05 1 9.901004556640303e-05 1 9.950984556640304e-05 1 9.951004556640304e-05 1 0.00010000984556640305 1 0.00010001004556640305 1 0.00010050984556640307 1 0.00010051004556640307 1 0.00010100984556640308 1 0.00010101004556640308 1 0.00010150984556640309 1 0.00010151004556640309 1 0.0001020098455664031 1 0.0001020100455664031 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00010771189158154771 1 0.00010771209158154771 1 0.0001082118915815477 1 0.0001082120915815477 1 0.00010871189158154768 1 0.00010871209158154768 1 0.00010921189158154767 1 0.00010921209158154767 1 0.00010971189158154765 1 0.00010971209158154765 1 0.00011021189158154764 1 0.00011021209158154764 1 0.00011071189158154762 1 0.00011071209158154762 1 0.00011121189158154761 1 0.00011121209158154761 1 0.00011171189158154759 1 0.00011171209158154759 1 0.00011221189158154758 1 0.00011221209158154758 1 0.00011241412374722472 1 0.00011241432374722472 1 0.0001179141237472247 1 0.0001179143237472247 1 0.00011841412374722469 1 0.00011841432374722469 1 0.00011891412374722467 1 0.00011891432374722467 1 0.00011941412374722466 1 0.00011941432374722466 1 0.00011991412374722464 1 0.00011991432374722464 1 0.00012041412374722463 1 0.00012041432374722463 1 0.00012091412374722461 1 0.00012091432374722461 1 0.00012141412374722461 1 0.00012141432374722461 1 0.00012191412374722461 1 0.00012191432374722461 1 0.0001224141237472246 1 0.00012241432374722458 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00012811667966227717 1 0.00012811687966227716 1 0.00012861667966227719 1 0.00012861687966227717 1 0.0001291166796622772 1 0.00012911687966227719 1 0.0001296166796622772 1 0.0001296168796622772 1 0.00013011667966227722 1 0.0001301168796622772 1 0.00013061667966227723 1 0.00013061687966227722 1 0.00013111667966227725 1 0.00013111687966227723 1 0.00013161667966227726 1 0.00013161687966227725 1 0.00013211667966227727 1 0.00013211687966227726 1 0.00013261667966227728 1 0.00013261687966227727 1 0.00013281929267817236 1 0.00013281949267817235 1 0.0001383192926781724 1 0.00013831949267817238 1 0.0001388192926781724 1 0.0001388194926781724 1 0.00013931929267817241 1 0.0001393194926781724 1 0.00013981929267817243 1 0.0001398194926781724 1 0.00014031929267817244 1 0.00014031949267817242 1 0.00014081929267817245 1 0.00014081949267817244 1 0.00014131929267817246 1 0.00014131949267817245 1 0.00014181929267817247 1 0.00014181949267817246 1 0.0001423192926781725 1 0.00014231949267817247 1 0.0001428192926781725 1 0.00014281949267817249 1 0.00014302214851901298 1 0.00014302234851901297 1 0.000148522148519013 1 0.000148522348519013 1 0.00014902214851901302 1 0.000149022348519013 1 0.00014952214851901303 1 0.00014952234851901302 1 0.00015002214851901304 1 0.00015002234851901303 1 0.00015052214851901305 1 0.00015052234851901304 1 0.00015102214851901307 1 0.00015102234851901305 1 0.00015152214851901308 1 0.00015152234851901306 1 0.0001520221485190131 1 0.00015202234851901308 1 0.0001525221485190131 1 0.0001525223485190131 1 0.00015302214851901311 1 0.0001530223485190131 1 0.00015322531083256498 1 0.00015322551083256497 1 0.000158725310832565 1 0.000158725510832565 1 0.00015922531083256502 1 0.000159225510832565 1 0.00015972531083256503 1 0.00015972551083256502 1 0.00016022531083256504 1 0.00016022551083256503 1 0.00016072531083256505 1 0.00016072551083256504 1 0.00016122531083256507 1 0.00016122551083256505 1 0.00016172531083256508 1 0.00016172551083256506 1 0.0001622253108325651 1 0.00016222551083256508 1 0.0001627253108325651 1 0.0001627255108325651 1 0.00016322531083256511 1 0.0001632255108325651 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001689286310398012 1 0.00016892883103980118 1 0.0001694286310398012 1 0.0001694288310398012 1 0.00016992863103980121 1 0.0001699288310398012 1 0.00017042863103980123 1 0.0001704288310398012 1 0.00017092863103980124 1 0.00017092883103980122 1 0.00017142863103980125 1 0.00017142883103980124 1 0.00017192863103980126 1 0.00017192883103980125 1 0.00017242863103980127 1 0.00017242883103980126 1 0.0001729286310398013 1 0.00017292883103980127 1 0.0001734286310398013 1 0.00017342883103980129 1 0.0001736321391540218 1 0.0001736323391540218 1 0.00017913213915402183 1 0.00017913233915402182 1 0.00017963213915402185 1 0.00017963233915402183 1 0.00018013213915402186 1 0.00018013233915402185 1 0.00018063213915402187 1 0.00018063233915402186 1 0.00018113213915402188 1 0.00018113233915402187 1 0.0001816321391540219 1 0.00018163233915402188 1 0.0001821321391540219 1 0.0001821323391540219 1 0.00018263213915402192 1 0.0001826323391540219 1 0.00018313213915402193 1 0.00018313233915402192 1 0.00018363213915402194 1 0.00018363233915402193 1 0.0001838358186013159 1 0.00018383601860131587 1 0.0001893358186013159 1 0.0001893360186013159 1 0.00018983581860131592 1 0.0001898360186013159 1 0.00019033581860131594 1 0.00019033601860131592 1 0.00019083581860131595 1 0.00019083601860131594 1 0.00019133581860131596 1 0.00019133601860131595 1 0.00019183581860131597 1 0.00019183601860131596 1 0.00019233581860131599 1 0.00019233601860131597 1 0.000192835818601316 1 0.00019283601860131598 1 0.000193335818601316 1 0.000193336018601316 1 0.00019383581860131602 1 0.000193836018601316 1 0.00019403971249211136 1 0.00019403991249211135 1 0.00019953971249211139 1 0.00019953991249211137 1 0.0002000397124921114 1 0.00020003991249211139 1 0.0002005397124921114 1 0.0002005399124921114 1 0.00020103971249211142 1 0.0002010399124921114 1 0.00020153971249211143 1 0.00020153991249211142 1 0.00020203971249211145 1 0.00020203991249211143 1 0.00020253971249211146 1 0.00020253991249211145 1 0.00020303971249211147 1 0.00020303991249211146 1 0.00020353971249211148 1 0.00020353991249211147 1 0.0002040397124921115 1 0.00020403991249211148 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00020974372730790412 1 0.0002097439273079041 1 0.00021024372730790413 1 0.00021024392730790412 1 0.00021074372730790414 1 0.00021074392730790413 1 0.00021124372730790415 1 0.00021124392730790414 1 0.00021174372730790416 1 0.00021174392730790415 1 0.00021224372730790418 1 0.00021224392730790416 1 0.0002127437273079042 1 0.00021274392730790418 1 0.0002132437273079042 1 0.0002132439273079042 1 0.0002137437273079042 1 0.0002137439273079042 1 0.00021424372730790423 1 0.0002142439273079042 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00021994808721675777 1 0.00021994828721675776 1 0.00022044808721675778 1 0.00022044828721675777 1 0.0002209480872167578 1 0.00022094828721675778 1 0.0002214480872167578 1 0.0002214482872167578 1 0.00022194808721675782 1 0.0002219482872167578 1 0.00022244808721675783 1 0.00022244828721675782 1 0.00022294808721675784 1 0.00022294828721675783 1 0.00022344808721675786 1 0.00022344828721675784 1 0.00022394808721675787 1 0.00022394828721675786 1 0.00022444808721675788 1 0.00022444828721675787 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023015261116331257 1 0.00023015281116331256 1 0.00023065261116331259 1 0.00023065281116331257 1 0.0002311526111633126 1 0.00023115281116331258 1 0.0002316526111633126 1 0.0002316528111633126 1 0.00023215261116331262 1 0.0002321528111633126 1 0.00023265261116331263 1 0.00023265281116331262 1 0.00023315261116331265 1 0.00023315281116331263 1 0.00023365261116331266 1 0.00023365281116331265 1 0.00023415261116331267 1 0.00023415281116331266 1 0.00023465261116331268 1 0.00023465281116331267 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024035725348777874 1 0.00024035745348777873 1 0.00024085725348777876 1 0.00024085745348777874 1 0.00024135725348777877 1 0.00024135745348777876 1 0.00024185725348777878 1 0.00024185745348777877 1 0.0002423572534877788 1 0.00024235745348777878 1 0.0002428572534877788 1 0.0002428574534877788 1 0.00024335725348777882 1 0.0002433574534877788 1 0.00024385725348777883 1 0.00024385745348777882 1 0.00024435725348777884 1 0.00024435745348777886 1 0.0002448572534877788 1 0.0002448574534877788 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025056213249421646 1 0.0002505623324942165 1 0.0002510621324942165 1 0.0002510623324942165 1 0.0002515621324942165 1 0.0002515623324942165 1 0.0002520621324942165 1 0.0002520623324942165 1 0.0002525621324942165 1 0.0002525623324942165 1 0.0002530621324942165 1 0.00025306233249421654 1 0.00025356213249421654 1 0.00025356233249421655 1 0.00025406213249421655 1 0.00025406233249421656 1 0.00025456213249421656 1 0.0002545623324942166 1 0.00025506213249421646 1 0.0002550623324942165 1 0.00025526732409400483 1 0.00025526752409400484 1 0.00026076732409400485 1 0.00026076752409400487 1 0.0002612673240940049 1 0.00026126752409400493 1 0.000261767324094005 1 0.000261767524094005 1 0.00026226732409400505 1 0.00026226752409400507 1 0.0002627673240940051 1 0.00026276752409400513 1 0.0002632673240940052 1 0.0002632675240940052 1 0.00026376732409400525 1 0.00026376752409400527 1 0.0002642673240940053 1 0.00026426752409400533 1 0.0002647673240940054 1 0.0002647675240940054 1 0.00026526732409400534 1 0.00026526752409400536 1 0.0002654725372742233 1 0.00026547273727422333 1 0.00027097253727422334 1 0.00027097273727422336 1 0.0002714725372742233 1 0.0002714727372742233 1 0.00027197253727422326 1 0.00027197273727422327 1 0.0002724725372742232 1 0.00027247273727422323 1 0.0002729725372742232 1 0.0002729727372742232 1 0.00027347253727422313 1 0.00027347273727422315 1 0.0002739725372742231 1 0.0002739727372742231 1 0.00027447253727422305 1 0.00027447273727422306 1 0.000274972537274223 1 0.000274972737274223 1 0.00027547253727422285 1 0.00027547273727422287 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002811781009094726 1 0.0002811783009094726 1 0.0002816781009094726 1 0.00028167830090947263 1 0.0002821781009094726 1 0.00028217830090947264 1 0.00028267810090947264 1 0.00028267830090947265 1 0.00028317810090947265 1 0.00028317830090947266 1 0.00028367810090947266 1 0.0002836783009094727 1 0.0002841781009094727 1 0.0002841783009094727 1 0.0002846781009094727 1 0.0002846783009094727 1 0.0002851781009094727 1 0.0002851783009094727 1 0.0002856781009094726 1 0.0002856783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.00029138383835494047 1 0.0002913840383549405 1 0.0002918838383549404 1 0.00029188403835494044 1 0.0002923838383549404 1 0.0002923840383549404 1 0.00029288383835494034 1 0.00029288403835494035 1 0.0002933838383549403 1 0.0002933840383549403 1 0.00029388383835494026 1 0.00029388403835494027 1 0.0002943838383549402 1 0.00029438403835494023 1 0.00029488383835494017 1 0.0002948840383549402 1 0.00029538383835494013 1 0.00029538403835494014 1 0.00029588383835494 1 0.00029588403835494 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003015896923277906 1 0.0003015898923277906 1 0.00030208969232779054 1 0.00030208989232779056 1 0.0003025896923277905 1 0.0003025898923277905 1 0.00030308969232779046 1 0.00030308989232779047 1 0.0003035896923277904 1 0.00030358989232779043 1 0.0003040896923277904 1 0.0003040898923277904 1 0.00030458969232779033 1 0.00030458989232779035 1 0.0003050896923277903 1 0.0003050898923277903 1 0.00030558969232779025 1 0.00030558989232779026 1 0.0003060896923277901 1 0.0003060898923277901 1 0.0003062957259554461 1 0.0003062959259554461 1 0.00031179572595544606 1 0.00031179592595544607 1 0.000312295725955446 1 0.00031229592595544603 1 0.000312795725955446 1 0.000312795925955446 1 0.00031329572595544593 1 0.00031329592595544595 1 0.0003137957259554459 1 0.0003137959259554459 1 0.00031429572595544585 1 0.00031429592595544586 1 0.0003147957259554458 1 0.0003147959259554458 1 0.00031529572595544576 1 0.0003152959259554458 1 0.0003157957259554457 1 0.00031579592595544574 1 0.00031629572595544557 1 0.0003162959259554456 1 0.0003165020377403174 1 0.0003165022377403174 1 0.00032200203774031743 1 0.00032200223774031745 1 0.0003225020377403175 1 0.0003225022377403175 1 0.00032300203774031757 1 0.0003230022377403176 1 0.00032350203774031763 1 0.00032350223774031765 1 0.0003240020377403177 1 0.0003240022377403177 1 0.00032450203774031777 1 0.0003245022377403178 1 0.00032500203774031783 1 0.00032500223774031785 1 0.0003255020377403179 1 0.0003255022377403179 1 0.00032600203774031796 1 0.000326002237740318 1 0.0003265020377403179 1 0.00032650223774031794 1 0.0003267084673472993 1 0.0003267086673472993 1 0.0003322084673472994 1 0.0003322086673472994 1 0.00033270846734729945 1 0.00033270866734729946 1 0.0003332084673472995 1 0.00033320866734729953 1 0.0003337084673472996 1 0.0003337086673472996 1 0.00033420846734729965 1 0.00033420866734729966 1 0.0003347084673472997 1 0.00033470866734729973 1 0.0003352084673472998 1 0.0003352086673472998 1 0.00033570846734729985 1 0.00033570866734729986 1 0.0003362084673472999 1 0.00033620866734729993 1 0.00033670846734729987 1 0.0003367086673472999 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034241523365255693 1 0.00034241543365255695 1 0.0003429152336525569 1 0.0003429154336525569 1 0.00034341523365255685 1 0.00034341543365255686 1 0.0003439152336525568 1 0.0003439154336525568 1 0.00034441523365255676 1 0.0003444154336525568 1 0.0003449152336525567 1 0.00034491543365255674 1 0.0003454152336525567 1 0.0003454154336525567 1 0.00034591523365255664 1 0.00034591543365255665 1 0.0003464152336525566 1 0.0003464154336525566 1 0.00034691523365255644 1 0.00034691543365255646 1 0.00034712205306404025 1 0.00034712225306404026 1 0.0003526220530640403 1 0.0003526222530640403 1 0.00035312205306404023 1 0.00035312225306404025 1 0.0003536220530640402 1 0.0003536222530640402 1 0.00035412205306404015 1 0.00035412225306404016 1 0.0003546220530640401 1 0.0003546222530640401 1 0.00035512205306404007 1 0.0003551222530640401 1 0.00035562205306404 1 0.00035562225306404004 1 0.00035612205306404 1 0.00035612225306404 1 0.00035662205306403994 1 0.00035662225306403995 1 0.0003571220530640398 1 0.0003571222530640398 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036282924646941807 1 0.0003628294464694181 1 0.0003633292464694181 1 0.0003633294464694181 1 0.0003638292464694181 1 0.0003638294464694181 1 0.0003643292464694181 1 0.0003643294464694181 1 0.0003648292464694181 1 0.00036482944646941813 1 0.00036532924646941813 1 0.00036532944646941814 1 0.00036582924646941814 1 0.00036582944646941815 1 0.00036632924646941815 1 0.00036632944646941817 1 0.00036682924646941817 1 0.0003668294464694182 1 0.00036732924646941807 1 0.0003673294464694181 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003730365334006625 1 0.0003730367334006625 1 0.0003735365334006625 1 0.0003735367334006625 1 0.0003740365334006625 1 0.00037403673340066253 1 0.0003745365334006625 1 0.00037453673340066254 1 0.00037503653340066254 1 0.00037503673340066255 1 0.00037553653340066255 1 0.00037553673340066256 1 0.00037603653340066256 1 0.0003760367334006626 1 0.0003765365334006626 1 0.0003765367334006626 1 0.0003770365334006626 1 0.0003770367334006626 1 0.0003775365334006625 1 0.0003775367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.0003832439556119043 1 0.0003832441556119043 1 0.00038374395561190425 1 0.00038374415561190427 1 0.0003842439556119042 1 0.0003842441556119042 1 0.00038474395561190417 1 0.0003847441556119042 1 0.0003852439556119041 1 0.00038524415561190414 1 0.0003857439556119041 1 0.0003857441556119041 1 0.00038624395561190404 1 0.00038624415561190406 1 0.000386743955611904 1 0.000386744155611904 1 0.00038724395561190396 1 0.00038724415561190397 1 0.0003877439556119038 1 0.0003877441556119038 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039345175422431377 1 0.0003934519542243138 1 0.0003939517542243138 1 0.0003939519542243138 1 0.0003944517542243138 1 0.0003944519542243138 1 0.0003949517542243138 1 0.0003949519542243138 1 0.0003954517542243138 1 0.00039545195422431383 1 0.0003959517542243138 1 0.00039595195422431384 1 0.00039645175422431384 1 0.00039645195422431385 1 0.00039695175422431385 1 0.00039695195422431386 1 0.00039745175422431386 1 0.0003974519542243139 1 0.00039795175422431377 1 0.0003979519542243138 1 0.00039815970887468034 1 0.00039815990887468036 1 0.0004036597088746804 1 0.00040365990887468044 1 0.0004041597088746805 1 0.0004041599088746805 1 0.00040465970887468056 1 0.00040465990887468057 1 0.0004051597088746806 1 0.00040515990887468064 1 0.0004056597088746807 1 0.0004056599088746807 1 0.00040615970887468076 1 0.00040615990887468077 1 0.0004066597088746808 1 0.00040665990887468084 1 0.0004071597088746809 1 0.0004071599088746809 1 0.00040765970887468095 1 0.00040765990887468097 1 0.0004081597088746809 1 0.0004081599088746809 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004138678210077549 1 0.0004138680210077549 1 0.00041436782100775496 1 0.00041436802100775497 1 0.000414867821007755 1 0.00041486802100775504 1 0.0004153678210077551 1 0.0004153680210077551 1 0.00041586782100775516 1 0.00041586802100775517 1 0.0004163678210077552 1 0.00041636802100775524 1 0.0004168678210077553 1 0.0004168680210077553 1 0.00041736782100775536 1 0.00041736802100775537 1 0.0004178678210077554 1 0.00041786802100775544 1 0.0004183678210077554 1 0.0004183680210077554 1 0.0004185760523824421 1 0.00041857625238244213 1 0.00042407605238244214 1 0.00042407625238244216 1 0.00042457605238244216 1 0.00042457625238244217 1 0.00042507605238244217 1 0.0004250762523824422 1 0.0004255760523824422 1 0.0004255762523824422 1 0.0004260760523824422 1 0.0004260762523824422 1 0.0004265760523824422 1 0.0004265762523824422 1 0.0004270760523824422 1 0.00042707625238244223 1 0.00042757605238244223 1 0.00042757625238244224 1 0.00042807605238244224 1 0.00042807625238244226 1 0.00042857605238244215 1 0.00042857625238244216 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043428458211686454 1 0.00043428478211686455 1 0.0004347845821168646 1 0.0004347847821168646 1 0.00043528458211686467 1 0.0004352847821168647 1 0.00043578458211686474 1 0.00043578478211686475 1 0.0004362845821168648 1 0.0004362847821168648 1 0.00043678458211686487 1 0.0004367847821168649 1 0.00043728458211686493 1 0.00043728478211686495 1 0.000437784582116865 1 0.000437784782116865 1 0.00043828458211686507 1 0.0004382847821168651 1 0.000438784582116865 1 0.00043878478211686504 1 0.00043899329473837736 1 0.00043899349473837737 1 0.0004444932947383774 1 0.0004444934947383774 1 0.0004449932947383774 1 0.0004449934947383774 1 0.0004454932947383774 1 0.0004454934947383774 1 0.0004459932947383774 1 0.00044599349473837743 1 0.00044649329473837743 1 0.00044649349473837745 1 0.00044699329473837744 1 0.00044699349473837746 1 0.00044749329473837746 1 0.00044749349473837747 1 0.00044799329473837747 1 0.0004479934947383775 1 0.0004484932947383775 1 0.0004484934947383775 1 0.0004489932947383774 1 0.0004489934947383774 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045470219161099484 1 0.00045470239161099485 1 0.0004552021916109948 1 0.0004552023916109948 1 0.00045570219161099475 1 0.00045570239161099477 1 0.0004562021916109947 1 0.0004562023916109947 1 0.00045670219161099467 1 0.0004567023916109947 1 0.0004572021916109946 1 0.00045720239161099464 1 0.0004577021916109946 1 0.0004577023916109946 1 0.00045820219161099454 1 0.00045820239161099456 1 0.0004587021916109945 1 0.0004587023916109945 1 0.00045920219161099435 1 0.00045920239161099436 1 0.00045941127816508494 1 0.00045941147816508496 1 0.00046491127816508497 1 0.000464911478165085 1 0.000465411278165085 1 0.000465411478165085 1 0.000465911278165085 1 0.000465911478165085 1 0.000466411278165085 1 0.000466411478165085 1 0.000466911278165085 1 0.00046691147816508503 1 0.00046741127816508503 1 0.00046741147816508504 1 0.00046791127816508504 1 0.00046791147816508506 1 0.00046841127816508505 1 0.00046841147816508507 1 0.00046891127816508507 1 0.0004689114781650851 1 0.00046941127816508497 1 0.000469411478165085 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004751205704165872 1 0.00047512077041658723 1 0.0004756205704165873 1 0.0004756207704165873 1 0.00047612057041658735 1 0.00047612077041658737 1 0.0004766205704165874 1 0.00047662077041658743 1 0.0004771205704165875 1 0.0004771207704165875 1 0.00047762057041658755 1 0.00047762077041658757 1 0.0004781205704165876 1 0.00047812077041658763 1 0.0004786205704165877 1 0.0004786207704165877 1 0.00047912057041658775 1 0.00047912077041658776 1 0.00047962057041658765 1 0.00047962077041658767 1 0.0004798301251576905 1 0.00047983032515769053 1 0.00048533012515769054 1 0.00048533032515769056 1 0.00048583012515769056 1 0.00048583032515769057 1 0.00048633012515769057 1 0.0004863303251576906 1 0.0004868301251576906 1 0.0004868303251576906 1 0.0004873301251576906 1 0.0004873303251576906 1 0.0004878301251576906 1 0.0004878303251576906 1 0.0004883301251576906 1 0.0004883303251576905 1 0.0004888301251576906 1 0.0004888303251576906 1 0.0004893301251576907 1 0.0004893303251576907 1 0.0004898301251576905 1 0.0004898303251576905 1 0.000490039780822236 1 0.000490039980822236 1 0.000495539780822236 1 0.000495539980822236 1 0.0004960397808222361 1 0.000496039980822236 1 0.0004965397808222361 1 0.0004965399808222361 1 0.0004970397808222362 1 0.0004970399808222362 1 0.0004975397808222363 1 0.0004975399808222362 1 0.0004980397808222363 1 0.0004980399808222363 1 0.0004985397808222364 1 0.0004985399808222364 1 0.0004990397808222365 1 0.0004990399808222364 1 0.0004995397808222365 1 0.0004995399808222365 1 0.0005000397808222364 1 0.0005000399808222363 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005057496159810823 1 0.0005057498159810823 1 0.0005062496159810824 1 0.0005062498159810824 1 0.0005067496159810825 1 0.0005067498159810824 1 0.0005072496159810825 1 0.0005072498159810825 1 0.0005077496159810826 1 0.0005077498159810826 1 0.0005082496159810827 1 0.0005082498159810826 1 0.0005087496159810827 1 0.0005087498159810827 1 0.0005092496159810828 1 0.0005092498159810828 1 0.0005097496159810829 1 0.0005097498159810828 1 0.0005102496159810827 1)
X8 __thm_sel_bld[0]_v thm_sel_bld[0] __thm_sel_bld[0]_s 0 inout_sw_mod
V9 __thm_sel_bld[0]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 0 1.0400399910590747e-05 0 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 1.2 5.1203456879677744e-05 1.2 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 0 0.00012261667966227715 0 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 0 0.00015322531083256498 0 0.00015322551083256497 0 0.0001634286310398012 0 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 0 0.00022465261116331255 0 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 1.2 0.0002858838383549405 1.2 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 0 0.0003062957259554461 0 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 0 0.00035732924646941804 0 0.00035732944646941806 1.2 0.00036753653340066246 1.2 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 1.2 0.00045941127816508494 1.2 0.00045941147816508496 1.2 0.0004696205704165872 1.2 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 0 0.0005002496159810823 0 0.0005002498159810822 0 0.0005102496159810827 0)
V10 __thm_sel_bld[0]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X11 __thm_sel_bld[1]_v thm_sel_bld[1] __thm_sel_bld[1]_s 0 inout_sw_mod
V12 __thm_sel_bld[1]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 1.2 0.00024506213249421644 1.2 0.00024506233249421645 1.2 0.00025526732409400483 1.2 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 0 0.0002756781009094726 0 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 0 0.0003165020377403174 0 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 0 0.00033691523365255696 0 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 0 0.00035732924646941804 0 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 1.2 0.00043899329473837736 1.2 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 1.2 0.00045941127816508494 1.2 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 1.2 0.000490039780822236 1.2 0.000490039980822236 0 0.0005002496159810823 0 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V13 __thm_sel_bld[1]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X14 __thm_sel_bld[2]_v thm_sel_bld[2] __thm_sel_bld[2]_s 0 inout_sw_mod
V15 __thm_sel_bld[2]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 1.2 2.0600911580126338e-05 1.2 2.060111158012634e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 0 4.1002390731437404e-05 0 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 0 0.00012261667966227715 0 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 1.2 0.00014302214851901298 1.2 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 0 0.0002042437273079041 0 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 0 0.0004287845821168645 0 0.0004287847821168645 1.2 0.00043899329473837736 1.2 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 0 0.0005102496159810827 0)
V16 __thm_sel_bld[2]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X17 __thm_sel_bld[3]_v thm_sel_bld[3] __thm_sel_bld[3]_s 0 inout_sw_mod
V18 __thm_sel_bld[3]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 0 0.00012261667966227715 0 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 1.2 0.00014302214851901298 1.2 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 1.2 0.0001736321391540218 1.2 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 0 0.00022465261116331255 0 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 1.2 0.0002654725372742233 1.2 0.00026547273727422333 0 0.0002756781009094726 0 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 0 0.0003062957259554461 0 0.0003062959259554461 0 0.0003165020377403174 0 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 0 0.00039815970887468034 0 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 0 0.0004185760523824421 0 0.00041857625238244213 0 0.0004287845821168645 0 0.0004287847821168645 1.2 0.00043899329473837736 1.2 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 1.2 0.00045941127816508494 1.2 0.00045941147816508496 1.2 0.0004696205704165872 1.2 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 0 0.0005002496159810823 0 0.0005002498159810822 0 0.0005102496159810827 0)
V19 __thm_sel_bld[3]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X20 __thm_sel_bld[4]_v thm_sel_bld[4] __thm_sel_bld[4]_s 0 inout_sw_mod
V21 __thm_sel_bld[4]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 0 1.0400399910590747e-05 0 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 1.2 5.1203456879677744e-05 1.2 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 0 0.00012261667966227715 0 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 1.2 0.00014302214851901298 1.2 0.00014302234851901297 0 0.00015322531083256498 0 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 1.2 0.0001736321391540218 1.2 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 0 0.0002042437273079041 0 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 0 0.00022465261116331255 0 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 1.2 0.00024506213249421644 1.2 0.00024506233249421645 1.2 0.00025526732409400483 1.2 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 0 0.0003062957259554461 0 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 0 0.00033691523365255696 0 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 0 0.00039815970887468034 0 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 0 0.0004287845821168645 0 0.0004287847821168645 1.2 0.00043899329473837736 1.2 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 1.2 0.00045941127816508494 1.2 0.00045941147816508496 1.2 0.0004696205704165872 1.2 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 0 0.0005002496159810823 0 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V22 __thm_sel_bld[4]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X23 __thm_sel_bld[5]_v thm_sel_bld[5] __thm_sel_bld[5]_s 0 inout_sw_mod
V24 __thm_sel_bld[5]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 1.2 5.1203456879677744e-05 1.2 5.1203656879677745e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 1.2 8.18080003149639e-05 1.2 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 0 0.00013281929267817236 0 0.00013281949267817235 1.2 0.00014302214851901298 1.2 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 0 0.0002042437273079041 0 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 0 0.0002756781009094726 0 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 0 0.0003165020377403174 0 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 0 0.0004185760523824421 0 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 1.2 0.00044920219161099487 1.2 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 1.2 0.0004696205704165872 1.2 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 0 0.0005102496159810827 0)
V25 __thm_sel_bld[5]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X26 __thm_sel_bld[6]_v thm_sel_bld[6] __thm_sel_bld[6]_s 0 inout_sw_mod
V27 __thm_sel_bld[6]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 0 1.0400399910590747e-05 0 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 0 4.1002390731437404e-05 0 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 0 0.00015322531083256498 0 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 1.2 0.00021444808721675775 1.2 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 1.2 0.0002654725372742233 1.2 0.00026547273727422333 0 0.0002756781009094726 0 0.0002756783009094726 1.2 0.0002858838383549405 1.2 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 0 0.00033691523365255696 0 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 0 0.00035732924646941804 0 0.00035732944646941806 1.2 0.00036753653340066246 1.2 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 0 0.0004287845821168645 0 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 1.2 0.00044920219161099487 1.2 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 1.2 0.0004696205704165872 1.2 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 1.2 0.000490039780822236 1.2 0.000490039980822236 0 0.0005002496159810823 0 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V28 __thm_sel_bld[6]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X29 __thm_sel_bld[7]_v thm_sel_bld[7] __thm_sel_bld[7]_s 0 inout_sw_mod
V30 __thm_sel_bld[7]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 0 1.0400399910590747e-05 0 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 0 0.00013281929267817236 0 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 1.2 0.00024506213249421644 1.2 0.00024506233249421645 1.2 0.00025526732409400483 1.2 0.00025526752409400484 1.2 0.0002654725372742233 1.2 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 0 0.00039815970887468034 0 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 0 0.0004185760523824421 0 0.00041857625238244213 0 0.0004287845821168645 0 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 1.2 0.00044920219161099487 1.2 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 1.2 0.0004696205704165872 1.2 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 1.2 0.000490039780822236 1.2 0.000490039980822236 0 0.0005002496159810823 0 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V31 __thm_sel_bld[7]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X32 __thm_sel_bld[8]_v thm_sel_bld[8] __thm_sel_bld[8]_s 0 inout_sw_mod
V33 __thm_sel_bld[8]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 0 0.00012261667966227715 0 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 1.2 0.00014302214851901298 1.2 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 0 0.0001634286310398012 0 0.00016342883103980118 1.2 0.0001736321391540218 1.2 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 1.2 0.00021444808721675775 1.2 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 1.2 0.00025526732409400483 1.2 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 0 0.0002756781009094726 0 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 0 0.0003062957259554461 0 0.0003062959259554461 0 0.0003165020377403174 0 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 0 0.00039815970887468034 0 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 0 0.0004185760523824421 0 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 1.2 0.00045941127816508494 1.2 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 1.2 0.000490039780822236 1.2 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 0 0.0005102496159810827 0)
V34 __thm_sel_bld[8]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X35 __thm_sel_bld[9]_v thm_sel_bld[9] __thm_sel_bld[9]_s 0 inout_sw_mod
V36 __thm_sel_bld[9]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 0 0.00013281929267817236 0 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 0 0.0001634286310398012 0 0.00016342883103980118 1.2 0.0001736321391540218 1.2 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 1.2 0.00025526732409400483 1.2 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 0 0.00033691523365255696 0 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 1.2 0.00036753653340066246 1.2 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 1.2 0.000490039780822236 1.2 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 0 0.0005102496159810827 0)
V37 __thm_sel_bld[9]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X38 __thm_sel_bld[10]_v thm_sel_bld[10] __thm_sel_bld[10]_s 0 inout_sw_mod
V39 __thm_sel_bld[10]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 0 4.1002390731437404e-05 0 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 0 0.00013281929267817236 0 0.00013281949267817235 1.2 0.00014302214851901298 1.2 0.00014302234851901297 0 0.00015322531083256498 0 0.00015322551083256497 0 0.0001634286310398012 0 0.00016342883103980118 1.2 0.0001736321391540218 1.2 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 1.2 0.0002654725372742233 1.2 0.00026547273727422333 0 0.0002756781009094726 0 0.0002756783009094726 1.2 0.0002858838383549405 1.2 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 0 0.0003062957259554461 0 0.0003062959259554461 0 0.0003165020377403174 0 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 0 0.00033691523365255696 0 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 1.2 0.00036753653340066246 1.2 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 0 0.0004185760523824421 0 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 1.2 0.00043899329473837736 1.2 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 1.2 0.00045941127816508494 1.2 0.00045941147816508496 1.2 0.0004696205704165872 1.2 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V40 __thm_sel_bld[10]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X41 __thm_sel_bld[11]_v thm_sel_bld[11] __thm_sel_bld[11]_s 0 inout_sw_mod
V42 __thm_sel_bld[11]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 1.2 2.0600911580126338e-05 1.2 2.060111158012634e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 0 4.1002390731437404e-05 0 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 0 8.18080003149639e-05 0 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 0 0.00015322531083256498 0 0.00015322551083256497 0 0.0001634286310398012 0 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 0 0.0002042437273079041 0 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 1.2 0.00024506213249421644 1.2 0.00024506233249421645 1.2 0.00025526732409400483 1.2 0.00025526752409400484 1.2 0.0002654725372742233 1.2 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 1.2 0.0002858838383549405 1.2 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 0 0.00039815970887468034 0 0.00039815990887468036 0 0.00040836782100775487 0 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V43 __thm_sel_bld[11]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X44 __thm_sel_bld[12]_v thm_sel_bld[12] __thm_sel_bld[12]_s 0 inout_sw_mod
V45 __thm_sel_bld[12]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 0 4.1002390731437404e-05 0 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 1.2 8.18080003149639e-05 1.2 8.18082003149639e-05 1.2 9.200984556640298e-05 1.2 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 0 0.00011241412374722472 0 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 0 0.0001634286310398012 0 0.00016342883103980118 1.2 0.0001736321391540218 1.2 0.0001736323391540218 0 0.0001838358186013159 0 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 0 0.0002042437273079041 0 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 1.2 0.00023485725348777872 1.2 0.0002348574534877787 1.2 0.00024506213249421644 1.2 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 1.2 0.0002654725372742233 1.2 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 1.2 0.00034712205306404025 1.2 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 1.2 0.00036753653340066246 1.2 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 0 0.0004287845821168645 0 0.0004287847821168645 1.2 0.00043899329473837736 1.2 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 0 0.0005102496159810827 0)
V46 __thm_sel_bld[12]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X47 __thm_sel_bld[13]_v thm_sel_bld[13] __thm_sel_bld[13]_s 0 inout_sw_mod
V48 __thm_sel_bld[13]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 0 1.0400399910590747e-05 0 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 0 4.1002390731437404e-05 0 4.1002590731437404e-05 0 5.1203456879677744e-05 0 5.1203656879677745e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 1.2 8.18080003149639e-05 1.2 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 1.2 0.00010221189158154771 1.2 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 0 0.00013281929267817236 0 0.00013281949267817235 1.2 0.00014302214851901298 1.2 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 1.2 0.0001736321391540218 1.2 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 0 0.0002042437273079041 0 0.00020424392730790408 1.2 0.00021444808721675775 1.2 0.00021444828721675773 1.2 0.00022465261116331255 1.2 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 1.2 0.0002654725372742233 1.2 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 1.2 0.0002960896923277906 1.2 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 1.2 0.0003267084673472993 1.2 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 0 0.0003777439556119043 0 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 0 0.00039815970887468034 0 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 0 0.0004185760523824421 0 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 0 0.0004798301251576905 0 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 0 0.0005102496159810827 0)
V49 __thm_sel_bld[13]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X50 __thm_sel_bld[14]_v thm_sel_bld[14] __thm_sel_bld[14]_s 0 inout_sw_mod
V51 __thm_sel_bld[14]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 1.2 1.0400399910590747e-05 1.2 1.0400599910590748e-05 0 2.0600911580126338e-05 0 2.060111158012634e-05 0 3.080158374751403e-05 0 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 1.2 5.1203456879677744e-05 1.2 5.1203656879677745e-05 0 6.140480297716098e-05 0 6.140500297716098e-05 0 7.160630340083568e-05 0 7.160650340083568e-05 1.2 8.18080003149639e-05 1.2 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 1.2 0.00012261667966227715 1.2 0.00012261687966227714 1.2 0.00013281929267817236 1.2 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 0 0.00015322531083256498 0 0.00015322551083256497 1.2 0.0001634286310398012 1.2 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 1.2 0.00019403971249211136 1.2 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 1.2 0.00021444808721675775 1.2 0.00021444828721675773 0 0.00022465261116331255 0 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 1.2 0.00024506213249421644 1.2 0.00024506233249421645 0 0.00025526732409400483 0 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 1.2 0.0002756781009094726 1.2 0.0002756783009094726 0 0.0002858838383549405 0 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 0 0.0003062957259554461 0 0.0003062959259554461 0 0.0003165020377403174 0 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 0 0.00036753653340066246 0 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 0 0.00038795175422431374 0 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 0 0.0004185760523824421 0 0.00041857625238244213 1.2 0.0004287845821168645 1.2 0.0004287847821168645 1.2 0.00043899329473837736 1.2 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 1.2 0.000490039780822236 1.2 0.000490039980822236 1.2 0.0005002496159810823 1.2 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V52 __thm_sel_bld[14]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
X53 __thm_sel_bld[15]_v thm_sel_bld[15] __thm_sel_bld[15]_s 0 inout_sw_mod
V54 __thm_sel_bld[15]_v 0 DC 0 PWL(0 0 2.001840282579421e-07 0 2.003840282579421e-07 0 1.0400399910590747e-05 0 1.0400599910590748e-05 1.2 2.0600911580126338e-05 1.2 2.060111158012634e-05 1.2 3.080158374751403e-05 1.2 3.080178374751403e-05 1.2 4.1002390731437404e-05 1.2 4.1002590731437404e-05 1.2 5.1203456879677744e-05 1.2 5.1203656879677745e-05 1.2 6.140480297716098e-05 1.2 6.140500297716098e-05 1.2 7.160630340083568e-05 1.2 7.160650340083568e-05 1.2 8.18080003149639e-05 1.2 8.18082003149639e-05 0 9.200984556640298e-05 0 9.201004556640298e-05 0 0.00010221189158154771 0 0.00010221209158154771 1.2 0.00011241412374722472 1.2 0.00011241432374722472 0 0.00012261667966227715 0 0.00012261687966227714 0 0.00013281929267817236 0 0.00013281949267817235 0 0.00014302214851901298 0 0.00014302234851901297 1.2 0.00015322531083256498 1.2 0.00015322551083256497 0 0.0001634286310398012 0 0.00016342883103980118 0 0.0001736321391540218 0 0.0001736323391540218 1.2 0.0001838358186013159 1.2 0.00018383601860131587 0 0.00019403971249211136 0 0.00019403991249211135 1.2 0.0002042437273079041 1.2 0.00020424392730790408 0 0.00021444808721675775 0 0.00021444828721675773 0 0.00022465261116331255 0 0.00022465281116331253 0 0.00023485725348777872 0 0.0002348574534877787 0 0.00024506213249421644 0 0.00024506233249421645 1.2 0.00025526732409400483 1.2 0.00025526752409400484 0 0.0002654725372742233 0 0.00026547273727422333 0 0.0002756781009094726 0 0.0002756783009094726 1.2 0.0002858838383549405 1.2 0.0002858840383549405 0 0.0002960896923277906 0 0.00029608989232779063 1.2 0.0003062957259554461 1.2 0.0003062959259554461 1.2 0.0003165020377403174 1.2 0.0003165022377403174 0 0.0003267084673472993 0 0.0003267086673472993 1.2 0.00033691523365255696 1.2 0.000336915433652557 0 0.00034712205306404025 0 0.00034712225306404026 1.2 0.00035732924646941804 1.2 0.00035732944646941806 1.2 0.00036753653340066246 1.2 0.0003675367334006625 1.2 0.0003777439556119043 1.2 0.00037774415561190434 1.2 0.00038795175422431374 1.2 0.00038795195422431375 1.2 0.00039815970887468034 1.2 0.00039815990887468036 1.2 0.00040836782100775487 1.2 0.0004083680210077549 1.2 0.0004185760523824421 1.2 0.00041857625238244213 0 0.0004287845821168645 0 0.0004287847821168645 0 0.00043899329473837736 0 0.00043899349473837737 0 0.00044920219161099487 0 0.0004492023916109949 0 0.00045941127816508494 0 0.00045941147816508496 0 0.0004696205704165872 0 0.0004696207704165872 1.2 0.0004798301251576905 1.2 0.00047983032515769053 0 0.000490039780822236 0 0.000490039980822236 0 0.0005002496159810823 0 0.0005002498159810822 1.2 0.0005102496159810827 1.2)
V55 __thm_sel_bld[15]_s 0 DC 1 PWL(0 1 2.001840282579421e-07 1 2.003840282579421e-07 1 1.0400399910590747e-05 1 1.0400599910590748e-05 1 2.0600911580126338e-05 1 2.060111158012634e-05 1 3.080158374751403e-05 1 3.080178374751403e-05 1 4.1002390731437404e-05 1 4.1002590731437404e-05 1 5.1203456879677744e-05 1 5.1203656879677745e-05 1 6.140480297716098e-05 1 6.140500297716098e-05 1 7.160630340083568e-05 1 7.160650340083568e-05 1 8.18080003149639e-05 1 8.18082003149639e-05 1 9.200984556640298e-05 1 9.201004556640298e-05 1 0.00010221189158154771 1 0.00010221209158154771 1 0.00011241412374722472 1 0.00011241432374722472 1 0.00012261667966227715 1 0.00012261687966227714 1 0.00013281929267817236 1 0.00013281949267817235 1 0.00014302214851901298 1 0.00014302234851901297 1 0.00015322531083256498 1 0.00015322551083256497 1 0.0001634286310398012 1 0.00016342883103980118 1 0.0001736321391540218 1 0.0001736323391540218 1 0.0001838358186013159 1 0.00018383601860131587 1 0.00019403971249211136 1 0.00019403991249211135 1 0.0002042437273079041 1 0.00020424392730790408 1 0.00021444808721675775 1 0.00021444828721675773 1 0.00022465261116331255 1 0.00022465281116331253 1 0.00023485725348777872 1 0.0002348574534877787 1 0.00024506213249421644 1 0.00024506233249421645 1 0.00025526732409400483 1 0.00025526752409400484 1 0.0002654725372742233 1 0.00026547273727422333 1 0.0002756781009094726 1 0.0002756783009094726 1 0.0002858838383549405 1 0.0002858840383549405 1 0.0002960896923277906 1 0.00029608989232779063 1 0.0003062957259554461 1 0.0003062959259554461 1 0.0003165020377403174 1 0.0003165022377403174 1 0.0003267084673472993 1 0.0003267086673472993 1 0.00033691523365255696 1 0.000336915433652557 1 0.00034712205306404025 1 0.00034712225306404026 1 0.00035732924646941804 1 0.00035732944646941806 1 0.00036753653340066246 1 0.0003675367334006625 1 0.0003777439556119043 1 0.00037774415561190434 1 0.00038795175422431374 1 0.00038795195422431375 1 0.00039815970887468034 1 0.00039815990887468036 1 0.00040836782100775487 1 0.0004083680210077549 1 0.0004185760523824421 1 0.00041857625238244213 1 0.0004287845821168645 1 0.0004287847821168645 1 0.00043899329473837736 1 0.00043899349473837737 1 0.00044920219161099487 1 0.0004492023916109949 1 0.00045941127816508494 1 0.00045941147816508496 1 0.0004696205704165872 1 0.0004696207704165872 1 0.0004798301251576905 1 0.00047983032515769053 1 0.000490039780822236 1 0.000490039980822236 1 0.0005002496159810823 1 0.0005002498159810822 1 0.0005102496159810827 1)
.probe ph_in[0] thm_sel_bld[0] ph_out thm_sel_bld[1] thm_sel_bld[2] ph_in[1]
.ic
.tran 5.102496159810827e-09 0.0005102496159810827
.end
